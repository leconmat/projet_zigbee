#  Last Change on: Thu Oct 21 13:18:13 2010
#  Owner: austriamicrosystems
#  Hit-Kit: Digital

#******
# Preview export LEF
#
#        Preview sub-version 5.10.41.500.6.138
#
# REF LIBS: IOLIB_4M
# TECH LIB NAME: TECH_C35B4
#******

VERSION 5.4 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 1000  ;
END UNITS

MANUFACTURINGGRID    0.025000 ;

SITE ioSite_P
    SYMMETRY Y  ;
    CLASS PAD  ;
    SIZE 100.000 BY 340.400 ;
END ioSite_P

SITE corner_P
    SYMMETRY R90  ;
    CLASS PAD  ;
    SIZE 340.400 BY 340.400 ;
END corner_P

MACRO GND3RP
    CLASS PAD ;
    FOREIGN GND3RP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
      #      CLASS CORE ;
        LAYER MET2 ;
        RECT  11.550 331.000 46.550 335.000 ;
        END
    END A
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 177.550 100.000 252.250 ;
        RECT  0.000 177.550 2.200 252.250 ;
        END
    END vdd3o!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 255.650 100.000 280.750 ;
        RECT  0.000 255.650 2.200 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 314.400 100.000 334.500 ;
        RECT  0.000 314.400 2.200 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 99.950 100.000 174.650 ;
        RECT  0.000 99.950 2.200 174.650 ;
        END
    END gnd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 282.550 100.000 312.650 ;
        RECT  0.000 282.550 2.200 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 330.200 ;
        RECT  0.000 -5.400 10.750 335.000 ;
        RECT  89.250 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  3.000 -5.400 97.000 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 335.000 ;
    END
END GND3RP

MACRO GND3OP
    CLASS PAD ;
    FOREIGN GND3OP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET4 ;
        RECT  5.500 3.050 94.850 92.000 ;
        END
    END A
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 177.550 100.000 252.250 ;
        RECT  0.000 177.550 2.200 252.250 ;
        END
    END vdd3o!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 255.650 100.000 280.750 ;
        RECT  0.000 255.650 2.200 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 314.400 100.000 334.500 ;
        RECT  0.000 314.400 2.200 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 99.950 100.000 174.650 ;
        RECT  0.000 99.950 2.200 174.650 ;
        END
    END gnd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 282.550 100.000 312.650 ;
        RECT  0.000 282.550 2.200 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  3.000 -5.400 97.000 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 2.250 ;
        RECT  0.000 -5.400 4.700 335.000 ;
        RECT  95.650 -5.400 97.500 335.000 ;
        RECT  0.000 92.800 100.000 335.000 ;
    END
END GND3OP

MACRO GND3IP
    CLASS PAD ;
    FOREIGN GND3IP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
            CLASS CORE ;
        LAYER MET2 ;
        RECT  11.550 331.000 46.550 335.000 ;
        END
    END A
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 177.550 100.000 252.250 ;
        RECT  0.000 177.550 2.200 252.250 ;
        END
    END vdd3o!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 255.650 100.000 280.750 ;
        RECT  0.000 255.650 2.200 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 314.400 100.000 334.500 ;
        RECT  0.000 314.400 2.200 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 99.950 100.000 174.650 ;
        RECT  0.000 99.950 2.200 174.650 ;
        END
    END gnd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 282.550 100.000 312.650 ;
        RECT  0.000 282.550 2.200 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 330.200 ;
        RECT  0.000 -5.400 10.750 335.000 ;
        RECT  89.250 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  3.000 -5.400 97.000 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 335.000 ;
    END
END GND3IP

MACRO GND3ALLP
    CLASS PAD ;
    FOREIGN GND3ALLP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
            CLASS CORE ;
        LAYER MET2 ;
        RECT  11.550 331.000 46.550 335.000 ;
        END
    END A
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 177.550 100.000 252.250 ;
        RECT  0.000 177.550 2.200 252.250 ;
        END
    END vdd3o!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 255.650 100.000 280.750 ;
        RECT  0.000 255.650 2.200 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 314.400 100.000 334.500 ;
        RECT  0.000 314.400 2.200 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  99.150 99.950 100.000 174.650 ;
        RECT  0.000 99.950 0.650 174.650 ;
        END
    END gnd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 282.550 100.000 312.650 ;
        RECT  0.000 282.550 2.200 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 330.200 ;
        RECT  0.000 -5.400 10.750 335.000 ;
        RECT  89.250 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  1.450 -5.400 98.350 176.750 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  3.000 -5.400 97.000 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 335.000 ;
    END
END GND3ALLP

MACRO VDD3RP
    CLASS PAD ;
    FOREIGN VDD3RP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET4 ;
        RECT  5.500 3.050 94.850 92.000 ;
        END
        PORT
      #      CLASS CORE ;
        LAYER MET2 ;
        RECT  11.600 331.450 46.600 335.000 ;
        END
    END A
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 177.550 100.000 252.250 ;
        RECT  0.000 177.550 2.200 252.250 ;
        END
    END vdd3o!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 255.650 100.000 280.750 ;
        RECT  0.000 255.650 2.200 280.750 ;
        END
    END vdd3r2!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 282.550 100.000 312.650 ;
        RECT  0.000 282.550 2.200 312.650 ;
        END
    END gnd3r!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 314.400 100.000 334.500 ;
        RECT  0.000 314.400 2.200 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 99.950 100.000 174.650 ;
        RECT  0.000 99.950 2.200 174.650 ;
        END
    END gnd3o!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 330.650 ;
        RECT  0.000 -5.400 10.800 335.000 ;
        RECT  89.300 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  3.000 -5.400 97.000 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 2.250 ;
        RECT  0.000 -5.400 4.700 335.000 ;
        RECT  95.650 -5.400 97.500 335.000 ;
        RECT  0.000 92.800 100.000 335.000 ;
    END
END VDD3RP

MACRO VDD3OP
    CLASS PAD ;
    FOREIGN VDD3OP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET4 ;
        RECT  5.500 3.050 94.850 92.000 ;
        END
    END A
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 177.550 100.000 252.250 ;
        RECT  0.000 177.550 2.200 252.250 ;
        END
    END vdd3o!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 255.650 100.000 280.750 ;
        RECT  0.000 255.650 2.200 280.750 ;
        END
    END vdd3r2!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 282.550 100.000 312.650 ;
        RECT  0.000 282.550 2.200 312.650 ;
        END
    END gnd3r!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 314.400 100.000 334.500 ;
        RECT  0.000 314.400 2.200 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 99.950 100.000 174.650 ;
        RECT  0.000 99.950 2.200 174.650 ;
        END
    END gnd3o!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  3.000 -5.400 97.000 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 2.250 ;
        RECT  0.000 -5.400 4.700 335.000 ;
        RECT  95.650 -5.400 97.500 335.000 ;
        RECT  0.000 92.800 100.000 335.000 ;
    END
END VDD3OP

MACRO VDD3IP
    CLASS PAD ;
    FOREIGN VDD3IP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET4 ;
        RECT  5.500 3.050 94.850 92.000 ;
        END
        PORT
            CLASS CORE ;
        LAYER MET2 ;
        RECT  11.600 331.000 46.600 335.000 ;
        END
    END A
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 177.550 100.000 252.250 ;
        RECT  0.000 177.550 2.200 252.250 ;
        END
    END vdd3o!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 255.650 100.000 280.750 ;
        RECT  0.000 255.650 2.200 280.750 ;
        END
    END vdd3r2!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 282.550 100.000 312.650 ;
        RECT  0.000 282.550 2.200 312.650 ;
        END
    END gnd3r!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 314.400 100.000 334.500 ;
        RECT  0.000 314.400 2.200 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 99.950 100.000 174.650 ;
        RECT  0.000 99.950 2.200 174.650 ;
        END
    END gnd3o!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 330.200 ;
        RECT  0.000 -5.400 10.800 335.000 ;
        RECT  89.300 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  3.000 -5.400 97.000 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 2.250 ;
        RECT  0.000 -5.400 4.700 335.000 ;
        RECT  95.650 -5.400 97.500 335.000 ;
        RECT  0.000 92.800 100.000 335.000 ;
    END
END VDD3IP

MACRO VDD3ALLP
    CLASS PAD ;
    FOREIGN VDD3ALLP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET4 ;
        RECT  5.500 3.050 94.850 92.000 ;
        END
        PORT
            CLASS CORE ;
        LAYER MET2 ;
        RECT  11.600 331.000 46.600 335.000 ;
        END
    END A
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 177.550 100.000 252.250 ;
        RECT  0.000 177.550 2.200 252.250 ;
        END
    END vdd3o!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 255.650 100.000 280.750 ;
        RECT  0.000 255.650 2.200 280.750 ;
        END
    END vdd3r2!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 282.550 100.000 312.650 ;
        RECT  0.000 282.550 2.200 312.650 ;
        END
    END gnd3r!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  97.800 314.400 100.000 334.500 ;
        RECT  0.000 314.400 2.200 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  97.800 99.950 100.000 174.650 ;
        RECT  0.000 99.950 2.200 174.650 ;
        END
    END gnd3o!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 330.200 ;
        RECT  0.000 -5.400 10.800 335.000 ;
        RECT  89.300 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  3.000 -5.400 97.000 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 2.250 ;
        RECT  0.000 -5.400 4.700 335.000 ;
        RECT  95.650 -5.400 97.500 335.000 ;
        RECT  0.000 92.800 100.000 335.000 ;
    END
END VDD3ALLP

MACRO RAILPROTP
    CLASS PAD ;
    FOREIGN RAILPROTP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 75.100 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  72.900 177.550 75.100 252.250 ;
        RECT  0.000 177.550 2.200 252.250 ;
        END
    END vdd3o!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  72.900 255.650 75.100 280.750 ;
        RECT  0.000 255.650 2.200 280.750 ;
        END
    END vdd3r2!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  72.900 282.550 75.100 312.650 ;
        RECT  0.000 282.550 2.200 312.650 ;
        END
    END gnd3r!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  72.900 314.400 75.100 334.500 ;
        RECT  0.000 314.400 2.200 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  72.900 99.950 75.100 174.650 ;
        RECT  0.000 99.950 2.200 174.650 ;
        END
    END gnd3o!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 75.100 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 75.100 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 75.100 99.150 ;
        RECT  0.000 175.450 75.100 176.750 ;
        RECT  0.000 253.050 75.100 254.850 ;
        RECT  0.000 281.550 75.100 281.750 ;
        RECT  0.000 313.450 75.100 313.600 ;
        RECT  3.000 -5.400 72.100 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 75.100 335.000 ;
    END
END RAILPROTP

MACRO PWRCUT_DIG_P_DX
    CLASS PAD ;
    FOREIGN PWRCUT_DIG_P_DX 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 50.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  46.000 99.950 50.000 174.650 ;
        RECT  0.000 99.950 4.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  46.000 255.650 50.000 280.750 ;
        RECT  0.000 255.650 4.000 280.750 ;
        END
    END vdd3r2!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  46.000 282.550 50.000 312.650 ;
        RECT  0.000 282.550 4.000 312.650 ;
        END
    END gnd3r!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  46.000 314.400 50.000 334.500 ;
        RECT  0.000 314.400 4.000 334.500 ;
        END
    END vdd3r1!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  46.000 177.550 50.000 252.250 ;
        RECT  0.000 177.550 4.000 252.250 ;
        END
    END vdd3o!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 50.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 50.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 50.000 99.150 ;
        RECT  0.000 175.450 50.000 176.750 ;
        RECT  0.000 253.050 50.000 254.850 ;
        RECT  0.000 281.550 50.000 281.750 ;
        RECT  0.000 313.450 50.000 313.600 ;
        RECT  4.800 -5.400 45.200 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 50.000 335.000 ;
    END
END PWRCUT_DIG_P_DX

MACRO CORNERP
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN CORNERP -5.4 -5.4 ;
    ORIGIN 5.400 5.400 ;
    SIZE 340.400 BY 340.400 ;
    SYMMETRY R90 ;
    SITE corner_P ;
    PIN gnd3o!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  331.000 99.950 335.000 174.650 ;
        RECT  99.950 331.000 174.650 335.000 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  331.000 177.550 335.000 252.250 ;
        RECT  177.550 331.000 252.250 335.000 ;
        END
    END vdd3o!
    PIN vdd3r2!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  331.000 255.650 335.000 280.750 ;
        RECT  255.650 331.000 280.750 335.000 ;
        END
    END vdd3r2!
    PIN gnd3r!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  331.000 282.550 335.000 312.650 ;
        RECT  282.550 331.000 312.650 335.000 ;
        END
    END gnd3r!
    PIN vdd3r1!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  331.000 314.400 335.000 334.500 ;
        RECT  314.400 331.000 334.500 335.000 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  -5.400 -5.400 335.000 335.000 ;
        LAYER MET2 ;
        RECT  -5.400 -5.400 335.000 335.000 ;
        LAYER MET3 ;
        RECT  -5.400 -5.400 335.000 99.150 ;
        RECT  -5.400 175.450 335.000 176.750 ;
        RECT  -5.400 253.050 335.000 254.850 ;
        RECT  -5.400 281.550 335.000 281.750 ;
        RECT  -5.400 313.450 335.000 313.600 ;
        RECT  -5.400 -5.400 330.200 330.200 ;
        RECT  -5.400 -5.400 99.150 335.000 ;
        RECT  175.450 -5.400 176.750 335.000 ;
        RECT  253.050 -5.400 254.850 335.000 ;
        RECT  281.550 -5.400 281.750 335.000 ;
        RECT  313.450 -5.400 313.600 335.000 ;
        LAYER MET4 ;
        RECT  -5.400 -5.400 335.000 335.000 ;
    END
END CORNERP

MACRO PERI_SPACER_5_P
    CLASS PAD SPACER ;
    FOREIGN PERI_SPACER_5_P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 5.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN gnd3o!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 99.950 5.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3r1!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 314.400 5.000 334.500 ;
        END
    END vdd3r1!
    PIN gnd3r!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 282.550 5.000 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 255.650 5.000 280.750 ;
        END
    END vdd3r2!
    PIN vdd3o!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 177.550 5.000 252.250 ;
        END
    END vdd3o!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 5.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 5.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 313.450 5.000 313.600 ;
        RECT  0.000 281.550 5.000 281.750 ;
        RECT  0.000 253.050 5.000 254.850 ;
        RECT  0.000 175.450 5.000 176.750 ;
        RECT  0.000 -5.400 5.000 99.150 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 5.000 335.000 ;
    END
END PERI_SPACER_5_P

MACRO PERI_SPACER_50_P
    CLASS PAD SPACER ;
    FOREIGN PERI_SPACER_50_P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 50.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  40.000 99.950 50.000 174.650 ;
        RECT  0.000 99.950 10.000 174.650 ;
        END
    END gnd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 282.550 50.000 312.650 ;
        END
    END gnd3r!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  40.000 177.550 50.000 252.250 ;
        RECT  0.000 177.550 10.000 252.250 ;
        END
    END vdd3o!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  29.950 314.400 50.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 255.650 50.000 280.750 ;
        END
    END vdd3r2!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 50.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 50.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 313.450 50.000 313.600 ;
        RECT  20.850 313.450 29.150 335.000 ;
        RECT  0.000 281.550 50.000 281.750 ;
        RECT  0.000 -5.400 50.000 99.150 ;
        RECT  0.000 175.450 50.000 176.750 ;
        RECT  10.800 -5.400 39.200 254.850 ;
        RECT  0.000 253.050 50.000 254.850 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 50.000 335.000 ;
    END
END PERI_SPACER_50_P

MACRO PERI_SPACER_2_P
    CLASS PAD SPACER ;
    FOREIGN PERI_SPACER_2_P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 2.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN gnd3o!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 99.950 2.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3r1!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 314.400 2.000 334.500 ;
        END
    END vdd3r1!
    PIN gnd3r!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 282.550 2.000 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 255.650 2.000 280.750 ;
        END
    END vdd3r2!
    PIN vdd3o!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 177.550 2.000 252.250 ;
        END
    END vdd3o!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 2.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 2.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 313.450 2.000 313.600 ;
        RECT  0.000 281.550 2.000 281.750 ;
        RECT  0.000 253.050 2.000 254.850 ;
        RECT  0.000 175.450 2.000 176.750 ;
        RECT  0.000 -5.400 2.000 99.150 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 2.000 335.000 ;
    END
END PERI_SPACER_2_P

MACRO PERI_SPACER_20_P
    CLASS PAD SPACER ;
    FOREIGN PERI_SPACER_20_P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 20.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 177.550 20.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 282.550 20.000 312.650 ;
        END
    END gnd3r!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 99.950 20.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 314.400 20.000 334.500 ;
        END
    END vdd3r1!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 255.650 20.000 280.750 ;
        END
    END vdd3r2!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 20.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 20.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 313.450 20.000 313.600 ;
        RECT  0.000 281.550 20.000 281.750 ;
        RECT  0.000 253.050 20.000 254.850 ;
        RECT  0.000 175.450 20.000 176.750 ;
        RECT  0.000 -5.400 20.000 99.150 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 20.000 335.000 ;
    END
END PERI_SPACER_20_P

MACRO PERI_SPACER_1_P
    CLASS PAD SPACER ;
    FOREIGN PERI_SPACER_1_P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 1.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN gnd3o!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 99.950 1.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3r1!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 314.400 1.000 334.500 ;
        END
    END vdd3r1!
    PIN gnd3r!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 282.550 1.000 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 255.650 1.000 280.750 ;
        END
    END vdd3r2!
    PIN vdd3o!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 177.550 1.000 252.250 ;
        END
    END vdd3o!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 1.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 1.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 313.450 1.000 313.600 ;
        RECT  0.000 281.550 1.000 281.750 ;
        RECT  0.000 253.050 1.000 254.850 ;
        RECT  0.000 175.450 1.000 176.750 ;
        RECT  0.000 -5.400 1.000 99.150 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 1.000 335.000 ;
    END
END PERI_SPACER_1_P

MACRO PERI_SPACER_10_P
    CLASS PAD SPACER ;
    FOREIGN PERI_SPACER_10_P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 10.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN gnd3o!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 99.950 10.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3r1!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 314.400 10.000 334.500 ;
        END
    END vdd3r1!
    PIN gnd3r!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 282.550 10.000 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 255.650 10.000 280.750 ;
        END
    END vdd3r2!
    PIN vdd3o!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 177.550 10.000 252.250 ;
        END
    END vdd3o!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 10.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 10.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 313.450 10.000 313.600 ;
        RECT  0.000 281.550 10.000 281.750 ;
        RECT  0.000 253.050 10.000 254.850 ;
        RECT  0.000 175.450 10.000 176.750 ;
        RECT  0.000 -5.400 10.000 99.150 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 10.000 335.000 ;
    END
END PERI_SPACER_10_P

MACRO PERI_SPACER_100_P
    CLASS PAD SPACER ;
    FOREIGN PERI_SPACER_100_P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 335.000 ;
    END
END PERI_SPACER_100_P

MACRO PERI_SPACER_01_P
    CLASS PAD SPACER ;
    FOREIGN PERI_SPACER_01_P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 0.100 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN gnd3o!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 99.950 0.100 174.650 ;
        END
    END gnd3o!
    PIN vdd3r1!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 314.400 0.100 334.500 ;
        END
    END vdd3r1!
    PIN gnd3r!
        DIRECTION FEEDTHRU ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 282.550 0.100 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 255.650 0.100 280.750 ;
        END
    END vdd3r2!
    PIN vdd3o!
        DIRECTION FEEDTHRU ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 177.550 0.100 252.250 ;
        END
    END vdd3o!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 0.100 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 0.100 335.000 ;
        LAYER MET3 ;
        RECT  0.000 313.450 0.100 313.600 ;
        RECT  0.000 281.550 0.100 281.750 ;
        RECT  0.000 253.050 0.100 254.850 ;
        RECT  0.000 175.450 0.100 176.750 ;
        RECT  0.000 -5.400 0.100 99.150 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 0.100 335.000 ;
    END
END PERI_SPACER_01_P

MACRO ITUP
    CLASS PAD ;
    FOREIGN ITUP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ITUP

MACRO ITP
    CLASS PAD ;
    FOREIGN ITP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ITP

MACRO ITDP
    CLASS PAD ;
    FOREIGN ITDP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ITDP

MACRO ITCK8P
    CLASS PAD ;
    FOREIGN ITCK8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 186.752  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  46.650 326.950 54.750 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 326.150 ;
        RECT  0.000 -5.400 45.850 335.000 ;
        RECT  55.550 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ITCK8P

MACRO ITCK4P
    CLASS PAD ;
    FOREIGN ITCK4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 135.296  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  48.850 330.950 52.950 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 330.150 ;
        RECT  0.000 -5.400 48.050 335.000 ;
        RECT  53.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ITCK4P

MACRO ITCK2P
    CLASS PAD ;
    FOREIGN ITCK2P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 108.160  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  49.650 332.550 52.150 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 331.750 ;
        RECT  0.000 -5.400 48.850 335.000 ;
        RECT  52.950 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ITCK2P

MACRO ITCK16P
    CLASS PAD ;
    FOREIGN ITCK16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 105.536  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  37.850 318.950 53.950 335.050 ;
        RECT  15.850 288.150 30.850 303.150 ;
        RECT  10.500 269.400 18.600 277.500 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 268.600 ;
        RECT  0.450 -5.400 9.800 335.000 ;
        RECT  10.300 278.000 11.200 335.000 ;
        RECT  19.400 -5.400 100.000 287.350 ;
        RECT  0.000 278.300 100.000 287.350 ;
        RECT  0.450 278.300 12.900 335.000 ;
        RECT  31.650 -5.400 100.000 318.150 ;
        RECT  0.000 303.950 37.050 335.000 ;
        RECT  54.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ITCK16P

MACRO ISUP
    CLASS PAD ;
    FOREIGN ISUP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 94.656  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  67.800 334.450 68.400 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 67.000 335.000 ;
        RECT  69.200 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ISUP

MACRO ISP
    CLASS PAD ;
    FOREIGN ISP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 94.656  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  67.800 334.450 68.400 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 67.000 335.000 ;
        RECT  69.200 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ISP

MACRO ISDP
    CLASS PAD ;
    FOREIGN ISDP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 94.656  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  67.800 334.450 68.400 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 67.000 335.000 ;
        RECT  69.200 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ISDP

MACRO ICUP
    CLASS PAD ;
    FOREIGN ICUP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ICUP

MACRO ICP
    CLASS PAD ;
    FOREIGN ICP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ICP

MACRO ICDP
    CLASS PAD ;
    FOREIGN ICDP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ICDP

MACRO ICCK8P
    CLASS PAD ;
    FOREIGN ICCK8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 186.752  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  46.650 326.950 54.750 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 326.150 ;
        RECT  0.000 -5.400 45.850 335.000 ;
        RECT  55.550 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ICCK8P

MACRO ICCK4P
    CLASS PAD ;
    FOREIGN ICCK4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 135.296  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  48.850 330.950 52.950 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 330.150 ;
        RECT  0.000 -5.400 48.050 335.000 ;
        RECT  53.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ICCK4P

MACRO ICCK2P
    CLASS PAD ;
    FOREIGN ICCK2P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 108.160  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  49.650 332.550 52.150 335.050 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 331.750 ;
        RECT  0.000 -5.400 48.850 335.000 ;
        RECT  52.950 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ICCK2P

MACRO ICCK16P
    CLASS PAD ;
    FOREIGN ICCK16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 105.344  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  37.850 318.950 53.950 335.050 ;
        RECT  16.000 288.150 31.000 303.150 ;
        RECT  10.500 269.400 18.600 277.500 ;
        END
    END Y
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 268.600 ;
        RECT  0.450 -5.400 9.800 335.000 ;
        RECT  10.300 278.000 11.200 335.000 ;
        RECT  19.400 -5.400 100.000 287.350 ;
        RECT  0.000 278.300 100.000 287.350 ;
        RECT  0.450 278.300 12.850 335.000 ;
        RECT  31.800 -5.400 100.000 318.150 ;
        RECT  0.000 303.950 37.050 335.000 ;
        RECT  54.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END ICCK16P

MACRO CBU2P
    CLASS PAD ;
    FOREIGN CBU2P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 40.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 62.656  LAYER MET2  ;
        ANTENNAGATEAREA 8.400  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  15.100 334.450 15.700 335.050 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 108.864  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  6.400 332.550 8.900 335.050 ;
        END
    END Y
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 255.650 40.000 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 314.400 40.000 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  35.000 99.950 40.000 174.650 ;
        RECT  0.000 99.950 5.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  35.000 177.550 40.000 252.250 ;
        RECT  0.000 177.550 5.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 282.550 40.000 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 40.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 40.000 331.750 ;
        RECT  9.700 -5.400 40.000 333.650 ;
        RECT  0.000 -5.400 5.600 335.000 ;
        RECT  9.700 -5.400 14.300 335.000 ;
        RECT  16.500 -5.400 40.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 313.450 40.000 313.600 ;
        RECT  0.000 281.550 40.000 281.750 ;
        RECT  0.000 -5.400 40.000 99.150 ;
        RECT  0.000 175.450 40.000 176.750 ;
        RECT  5.800 -5.400 34.200 254.850 ;
        RECT  0.000 253.050 40.000 254.850 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 40.000 335.000 ;
    END
END CBU2P

MACRO CBU1P
    CLASS PAD ;
    FOREIGN CBU1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 40.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.008  LAYER MET2  ;
        ANTENNAGATEAREA 4.200  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  15.100 334.450 15.700 335.050 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 108.864  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  6.400 332.550 8.900 335.050 ;
        END
    END Y
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 255.650 40.000 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  0.000 314.400 40.000 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  35.000 99.950 40.000 174.650 ;
        RECT  0.000 99.950 5.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  35.000 177.550 40.000 252.250 ;
        RECT  0.000 177.550 5.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  0.000 282.550 40.000 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 40.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 40.000 331.750 ;
        RECT  9.700 -5.400 40.000 333.650 ;
        RECT  0.000 -5.400 5.600 335.000 ;
        RECT  9.700 -5.400 14.300 335.000 ;
        RECT  16.500 -5.400 40.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 313.450 40.000 313.600 ;
        RECT  0.000 281.550 40.000 281.750 ;
        RECT  0.000 -5.400 40.000 99.150 ;
        RECT  0.000 175.450 40.000 176.750 ;
        RECT  5.800 -5.400 34.200 254.850 ;
        RECT  0.000 253.050 40.000 254.850 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 40.000 335.000 ;
    END
END CBU1P

MACRO BUDU8P
    CLASS PAD ;
    FOREIGN BUDU8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDU8P

MACRO BUDU4P
    CLASS PAD ;
    FOREIGN BUDU4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDU4P

MACRO BUDU2P
    CLASS PAD ;
    FOREIGN BUDU2P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDU2P

MACRO BUDU24P
    CLASS PAD ;
    FOREIGN BUDU24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDU24P

MACRO BUDU1P
    CLASS PAD ;
    FOREIGN BUDU1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDU1P

MACRO BUDU16P
    CLASS PAD ;
    FOREIGN BUDU16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDU16P

MACRO BUDU12P
    CLASS PAD ;
    FOREIGN BUDU12P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDU12P

MACRO BUDD8P
    CLASS PAD ;
    FOREIGN BUDD8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDD8P

MACRO BUDD4P
    CLASS PAD ;
    FOREIGN BUDD4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDD4P

MACRO BUDD2P
    CLASS PAD ;
    FOREIGN BUDD2P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDD2P

MACRO BUDD24P
    CLASS PAD ;
    FOREIGN BUDD24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDD24P

MACRO BUDD1P
    CLASS PAD ;
    FOREIGN BUDD1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDD1P

MACRO BUDD16P
    CLASS PAD ;
    FOREIGN BUDD16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDD16P

MACRO BUDD12P
    CLASS PAD ;
    FOREIGN BUDD12P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BUDD12P

MACRO BU8SP
    CLASS PAD ;
    FOREIGN BU8SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU8SP

MACRO BU8SMP
    CLASS PAD ;
    FOREIGN BU8SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU8SMP

MACRO BU8P
    CLASS PAD ;
    FOREIGN BU8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU8P

MACRO BU4SMP
    CLASS PAD ;
    FOREIGN BU4SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU4SMP

MACRO BU4P
    CLASS PAD ;
    FOREIGN BU4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU4P

MACRO BU2P
    CLASS PAD ;
    FOREIGN BU2P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU2P

MACRO BU24SP
    CLASS PAD ;
    FOREIGN BU24SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU24SP

MACRO BU24SMP
    CLASS PAD ;
    FOREIGN BU24SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU24SMP

MACRO BU24P
    CLASS PAD ;
    FOREIGN BU24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU24P

MACRO BU1P
    CLASS PAD ;
    FOREIGN BU1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU1P

MACRO BU16SP
    CLASS PAD ;
    FOREIGN BU16SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU16SP

MACRO BU16SMP
    CLASS PAD ;
    FOREIGN BU16SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU16SMP

MACRO BU16P
    CLASS PAD ;
    FOREIGN BU16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU16P

MACRO BU12SP
    CLASS PAD ;
    FOREIGN BU12SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU12SP

MACRO BU12SMP
    CLASS PAD ;
    FOREIGN BU12SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU12SMP

MACRO BU12P
    CLASS PAD ;
    FOREIGN BU12P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.920  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  2.700 334.450 3.300 335.050 ;
        END
    END A
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 1.900 335.000 ;
        RECT  4.100 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BU12P

MACRO BT8SP
    CLASS PAD ;
    FOREIGN BT8SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT8SP

MACRO BT8SMP
    CLASS PAD ;
    FOREIGN BT8SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT8SMP

MACRO BT8P
    CLASS PAD ;
    FOREIGN BT8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT8P

MACRO BT4SMP
    CLASS PAD ;
    FOREIGN BT4SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT4SMP

MACRO BT4P
    CLASS PAD ;
    FOREIGN BT4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT4P

MACRO BT2P
    CLASS PAD ;
    FOREIGN BT2P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT2P

MACRO BT24SP
    CLASS PAD ;
    FOREIGN BT24SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT24SP

MACRO BT24SMP
    CLASS PAD ;
    FOREIGN BT24SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT24SMP

MACRO BT24P
    CLASS PAD ;
    FOREIGN BT24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT24P

MACRO BT1P
    CLASS PAD ;
    FOREIGN BT1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT1P

MACRO BT16SP
    CLASS PAD ;
    FOREIGN BT16SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT16SP

MACRO BT16SMP
    CLASS PAD ;
    FOREIGN BT16SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT16SMP

MACRO BT16P
    CLASS PAD ;
    FOREIGN BT16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT16P

MACRO BT12SP
    CLASS PAD ;
    FOREIGN BT12SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT12SP

MACRO BT12SMP
    CLASS PAD ;
    FOREIGN BT12SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT12SMP

MACRO BT12P
    CLASS PAD ;
    FOREIGN BT12P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BT12P

MACRO BBTU8SP
    CLASS PAD ;
    FOREIGN BBTU8SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU8SP

MACRO BBTU8SMP
    CLASS PAD ;
    FOREIGN BBTU8SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU8SMP

MACRO BBTU8P
    CLASS PAD ;
    FOREIGN BBTU8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU8P

MACRO BBTU4SMP
    CLASS PAD ;
    FOREIGN BBTU4SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU4SMP

MACRO BBTU4P
    CLASS PAD ;
    FOREIGN BBTU4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU4P

MACRO BBTU24SP
    CLASS PAD ;
    FOREIGN BBTU24SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU24SP

MACRO BBTU24SMP
    CLASS PAD ;
    FOREIGN BBTU24SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU24SMP

MACRO BBTU24P
    CLASS PAD ;
    FOREIGN BBTU24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU24P

MACRO BBTU1P
    CLASS PAD ;
    FOREIGN BBTU1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU1P

MACRO BBTU16SP
    CLASS PAD ;
    FOREIGN BBTU16SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU16SP

MACRO BBTU16SMP
    CLASS PAD ;
    FOREIGN BBTU16SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU16SMP

MACRO BBTU16P
    CLASS PAD ;
    FOREIGN BBTU16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTU16P

MACRO BBTD8SP
    CLASS PAD ;
    FOREIGN BBTD8SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD8SP

MACRO BBTD8SMP
    CLASS PAD ;
    FOREIGN BBTD8SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD8SMP

MACRO BBTD8P
    CLASS PAD ;
    FOREIGN BBTD8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD8P

MACRO BBTD4SMP
    CLASS PAD ;
    FOREIGN BBTD4SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD4SMP

MACRO BBTD4P
    CLASS PAD ;
    FOREIGN BBTD4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD4P

MACRO BBTD24SP
    CLASS PAD ;
    FOREIGN BBTD24SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD24SP

MACRO BBTD24SMP
    CLASS PAD ;
    FOREIGN BBTD24SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD24SMP

MACRO BBTD24P
    CLASS PAD ;
    FOREIGN BBTD24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD24P

MACRO BBTD1P
    CLASS PAD ;
    FOREIGN BBTD1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD1P

MACRO BBTD16SP
    CLASS PAD ;
    FOREIGN BBTD16SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD16SP

MACRO BBTD16SMP
    CLASS PAD ;
    FOREIGN BBTD16SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD16SMP

MACRO BBTD16P
    CLASS PAD ;
    FOREIGN BBTD16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBTD16P

MACRO BBT8SP
    CLASS PAD ;
    FOREIGN BBT8SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT8SP

MACRO BBT8SMP
    CLASS PAD ;
    FOREIGN BBT8SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT8SMP

MACRO BBT8P
    CLASS PAD ;
    FOREIGN BBT8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT8P

MACRO BBT4SMP
    CLASS PAD ;
    FOREIGN BBT4SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT4SMP

MACRO BBT4P
    CLASS PAD ;
    FOREIGN BBT4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT4P

MACRO BBT24SP
    CLASS PAD ;
    FOREIGN BBT24SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT24SP

MACRO BBT24SMP
    CLASS PAD ;
    FOREIGN BBT24SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT24SMP

MACRO BBT24P
    CLASS PAD ;
    FOREIGN BBT24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT24P

MACRO BBT1P
    CLASS PAD ;
    FOREIGN BBT1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT1P

MACRO BBT16SP
    CLASS PAD ;
    FOREIGN BBT16SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT16SP

MACRO BBT16SMP
    CLASS PAD ;
    FOREIGN BBT16SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT16SMP

MACRO BBT16P
    CLASS PAD ;
    FOREIGN BBT16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 63.936  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBT16P

MACRO BBSU8SP
    CLASS PAD ;
    FOREIGN BBSU8SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU8SP

MACRO BBSU8SMP
    CLASS PAD ;
    FOREIGN BBSU8SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU8SMP

MACRO BBSU8P
    CLASS PAD ;
    FOREIGN BBSU8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU8P

MACRO BBSU4SMP
    CLASS PAD ;
    FOREIGN BBSU4SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU4SMP

MACRO BBSU4P
    CLASS PAD ;
    FOREIGN BBSU4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU4P

MACRO BBSU24SP
    CLASS PAD ;
    FOREIGN BBSU24SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU24SP

MACRO BBSU24SMP
    CLASS PAD ;
    FOREIGN BBSU24SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU24SMP

MACRO BBSU24P
    CLASS PAD ;
    FOREIGN BBSU24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU24P

MACRO BBSU1P
    CLASS PAD ;
    FOREIGN BBSU1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU1P

MACRO BBSU16SP
    CLASS PAD ;
    FOREIGN BBSU16SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU16SP

MACRO BBSU16SMP
    CLASS PAD ;
    FOREIGN BBSU16SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU16SMP

MACRO BBSU16P
    CLASS PAD ;
    FOREIGN BBSU16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSU16P

MACRO BBSD8SP
    CLASS PAD ;
    FOREIGN BBSD8SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD8SP

MACRO BBSD8SMP
    CLASS PAD ;
    FOREIGN BBSD8SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD8SMP

MACRO BBSD8P
    CLASS PAD ;
    FOREIGN BBSD8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD8P

MACRO BBSD4SMP
    CLASS PAD ;
    FOREIGN BBSD4SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD4SMP

MACRO BBSD4P
    CLASS PAD ;
    FOREIGN BBSD4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD4P

MACRO BBSD24SP
    CLASS PAD ;
    FOREIGN BBSD24SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD24SP

MACRO BBSD24SMP
    CLASS PAD ;
    FOREIGN BBSD24SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD24SMP

MACRO BBSD24P
    CLASS PAD ;
    FOREIGN BBSD24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD24P

MACRO BBSD1P
    CLASS PAD ;
    FOREIGN BBSD1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD1P

MACRO BBSD16SP
    CLASS PAD ;
    FOREIGN BBSD16SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD16SP

MACRO BBSD16SMP
    CLASS PAD ;
    FOREIGN BBSD16SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD16SMP

MACRO BBSD16P
    CLASS PAD ;
    FOREIGN BBSD16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBSD16P

MACRO BBS8SP
    CLASS PAD ;
    FOREIGN BBS8SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS8SP

MACRO BBS8SMP
    CLASS PAD ;
    FOREIGN BBS8SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS8SMP

MACRO BBS8P
    CLASS PAD ;
    FOREIGN BBS8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS8P

MACRO BBS4SMP
    CLASS PAD ;
    FOREIGN BBS4SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS4SMP

MACRO BBS4P
    CLASS PAD ;
    FOREIGN BBS4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS4P

MACRO BBS24SP
    CLASS PAD ;
    FOREIGN BBS24SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS24SP

MACRO BBS24SMP
    CLASS PAD ;
    FOREIGN BBS24SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS24SMP

MACRO BBS24P
    CLASS PAD ;
    FOREIGN BBS24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS24P

MACRO BBS1P
    CLASS PAD ;
    FOREIGN BBS1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS1P

MACRO BBS16SP
    CLASS PAD ;
    FOREIGN BBS16SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS16SP

MACRO BBS16SMP
    CLASS PAD ;
    FOREIGN BBS16SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS16SMP

MACRO BBS16P
    CLASS PAD ;
    FOREIGN BBS16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.152  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.450 4.900 335.050 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 104.256  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.450 75.900 335.050 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.512  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.450 10.950 335.050 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  74.500 282.550 75.300 313.000 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.650 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 73.700 313.600 ;
        RECT  76.100 313.450 100.000 313.600 ;
        RECT  20.850 314.400 79.150 334.500 ;
        RECT  20.850 313.450 73.700 335.000 ;
        RECT  76.100 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBS16P

MACRO BBCU8SP
    CLASS PAD ;
    FOREIGN BBCU8SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU8SP

MACRO BBCU8SMP
    CLASS PAD ;
    FOREIGN BBCU8SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU8SMP

MACRO BBCU8P
    CLASS PAD ;
    FOREIGN BBCU8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU8P

MACRO BBCU4SMP
    CLASS PAD ;
    FOREIGN BBCU4SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU4SMP

MACRO BBCU4P
    CLASS PAD ;
    FOREIGN BBCU4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU4P

MACRO BBCU24SP
    CLASS PAD ;
    FOREIGN BBCU24SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU24SP

MACRO BBCU24SMP
    CLASS PAD ;
    FOREIGN BBCU24SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU24SMP

MACRO BBCU24P
    CLASS PAD ;
    FOREIGN BBCU24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU24P

MACRO BBCU1P
    CLASS PAD ;
    FOREIGN BBCU1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU1P

MACRO BBCU16SP
    CLASS PAD ;
    FOREIGN BBCU16SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU16SP

MACRO BBCU16SMP
    CLASS PAD ;
    FOREIGN BBCU16SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU16SMP

MACRO BBCU16P
    CLASS PAD ;
    FOREIGN BBCU16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCU16P

MACRO BBCD8SP
    CLASS PAD ;
    FOREIGN BBCD8SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD8SP

MACRO BBCD8SMP
    CLASS PAD ;
    FOREIGN BBCD8SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD8SMP

MACRO BBCD8P
    CLASS PAD ;
    FOREIGN BBCD8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD8P

MACRO BBCD4SMP
    CLASS PAD ;
    FOREIGN BBCD4SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD4SMP

MACRO BBCD4P
    CLASS PAD ;
    FOREIGN BBCD4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD4P

MACRO BBCD24SP
    CLASS PAD ;
    FOREIGN BBCD24SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD24SP

MACRO BBCD24SMP
    CLASS PAD ;
    FOREIGN BBCD24SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD24SMP

MACRO BBCD24P
    CLASS PAD ;
    FOREIGN BBCD24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD24P

MACRO BBCD1P
    CLASS PAD ;
    FOREIGN BBCD1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD1P

MACRO BBCD16SP
    CLASS PAD ;
    FOREIGN BBCD16SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD16SP

MACRO BBCD16SMP
    CLASS PAD ;
    FOREIGN BBCD16SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD16SMP

MACRO BBCD16P
    CLASS PAD ;
    FOREIGN BBCD16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBCD16P

MACRO BBC8SP
    CLASS PAD ;
    FOREIGN BBC8SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC8SP

MACRO BBC8SMP
    CLASS PAD ;
    FOREIGN BBC8SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC8SMP

MACRO BBC8P
    CLASS PAD ;
    FOREIGN BBC8P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC8P

MACRO BBC4SMP
    CLASS PAD ;
    FOREIGN BBC4SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC4SMP

MACRO BBC4P
    CLASS PAD ;
    FOREIGN BBC4P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC4P

MACRO BBC24SP
    CLASS PAD ;
    FOREIGN BBC24SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC24SP

MACRO BBC24SMP
    CLASS PAD ;
    FOREIGN BBC24SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC24SMP

MACRO BBC24P
    CLASS PAD ;
    FOREIGN BBC24P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC24P

MACRO BBC1P
    CLASS PAD ;
    FOREIGN BBC1P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 2.800  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC1P

MACRO BBC16SP
    CLASS PAD ;
    FOREIGN BBC16SP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC16SP

MACRO BBC16SMP
    CLASS PAD ;
    FOREIGN BBC16SMP 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC16SMP

MACRO BBC16P
    CLASS PAD ;
    FOREIGN BBC16P 0 -5.4 ;
    ORIGIN 0.000 5.400 ;
    SIZE 100.000 BY 340.400 ;
    SYMMETRY R90 ;
    SITE ioSite_P ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER MET4 ;
        RECT  2.500 0.000 97.500 95.000 ;
        END
    END PAD
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 73.088  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  4.300 334.400 4.900 335.000 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 93.760  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  75.300 334.400 75.900 335.000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 72.448  LAYER MET2  ;
        ANTENNAGATEAREA 5.600  LAYER MET2  ;
        PORT
        LAYER MET2 ;
        RECT  10.350 334.400 10.950 335.000 ;
        END
    END A
    PIN gnd3o!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  85.000 99.950 100.000 174.650 ;
        RECT  0.000 99.950 15.000 174.650 ;
        END
    END gnd3o!
    PIN vdd3o!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  85.000 177.550 100.000 252.250 ;
        RECT  0.000 177.550 15.000 252.250 ;
        END
    END vdd3o!
    PIN gnd3r!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER MET3 ;
        RECT  69.950 282.550 100.000 312.650 ;
        RECT  0.000 282.550 30.050 312.650 ;
        END
    END gnd3r!
    PIN vdd3r2!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  74.950 255.650 100.000 280.750 ;
        RECT  0.000 255.650 25.050 280.750 ;
        END
    END vdd3r2!
    PIN vdd3r1!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER MET3 ;
        RECT  79.950 314.400 100.000 334.500 ;
        RECT  0.000 314.400 20.050 334.500 ;
        END
    END vdd3r1!
    OBS
        LAYER MET1 ;
        RECT  0.000 -5.400 100.000 335.000 ;
        LAYER MET2 ;
        RECT  0.000 -5.400 100.000 333.600 ;
        RECT  0.000 -5.400 3.500 335.000 ;
        RECT  5.700 -5.400 9.550 335.000 ;
        RECT  11.750 -5.400 74.500 335.000 ;
        RECT  76.700 -5.400 100.000 335.000 ;
        LAYER MET3 ;
        RECT  0.000 -5.400 100.000 99.150 ;
        RECT  0.000 175.450 100.000 176.750 ;
        RECT  15.800 -5.400 84.200 254.850 ;
        RECT  0.000 253.050 100.000 254.850 ;
        RECT  25.850 -5.400 74.150 281.750 ;
        RECT  0.000 281.550 100.000 281.750 ;
        RECT  30.850 -5.400 69.150 335.000 ;
        RECT  0.000 313.450 100.000 313.600 ;
        RECT  20.850 313.450 79.150 335.000 ;
        LAYER MET4 ;
        RECT  0.000 -5.400 100.000 -0.800 ;
        RECT  0.000 -5.400 1.700 335.000 ;
        RECT  0.000 95.800 100.000 335.000 ;
    END
END BBC16P

END LIBRARY
