module fifo_rx				
#(
					parameter WIDTH = 8,
					parameter DEPTH = 64
)		
(
					input logic clk, // horloge systeme 
					input logic reset_n,
					input logic en_cdr,
					// APB signals
					input logic data_in,
					input logic psel,
					input logic pwrite,
					input logic penable,
					output logic pready,
					output logic pslverr,
					// Output Tx
					output logic [WIDTH-1:0] prdata, 
					output reg mem_state // 0 memoire vide, 1 memoire remplie ou partiellement remplie
);


//////////////////////////////////////////////
//////////// Internal signals
//////////////////////////////////////////////
// Memory signals 
parameter PTR_WIDTH = $clog2(DEPTH);
logic [WIDTH-1:0] mem [DEPTH-1:0];
// Memory pointers	
logic [PTR_WIDTH:0] wr_ptr, rd_ptr;
// Memory flag
logic full;  
logic empty; 
reg [7:0] shift_register;
reg [WIDTH-1:0] i = 0;
reg en_cdr_prec;
assign pready = 1'b1;



/////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////// BEGIN MEMORY LOGIC ////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////

always_comb begin
	if((wr_ptr[PTR_WIDTH-1:0]) == (rd_ptr[PTR_WIDTH-1:0])) begin
		full = (wr_ptr[PTR_WIDTH]) ^ (rd_ptr[PTR_WIDTH]); // carry different => full 
		empty = wr_ptr[PTR_WIDTH] ~^ rd_ptr[PTR_WIDTH]; // carry identique => empty
	end
	else begin
		full = 0;
		empty = 0;
	end
end

// Memory state logic 
always_comb begin 
	if (full == 1'b1) begin
		mem_state = 1'b0; // Memoire vide 
	end
	else
		mem_state = 1'b1;
end

// APB Error logic
always_comb begin
	if (empty == 1) begin 
		pslverr = 1'b1; // Memoire pleine 
	end
	else 
		pslverr = 1'b0;
end

/////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////// END MEMORY LOGIC //////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////


/////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////// BEGIN WRITE LOGIC /////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////

assign wr_en = !en_cdr_prec && en_cdr && !full ;

// Shift register SERIAL IN PARALLEL OUT 
always @(posedge clk, negedge reset_n) begin
	if (!reset_n) begin
		shift_register <= 8'b00000000;
	end
	else begin
		if (i >= WIDTH)
			i <= 0;
		else begin
			shift_register[i] <= data_in;
			i <= i + 1;
		end
	end
end

always_ff @(posedge clk, negedge reset_n) begin
	if(~reset_n) begin
		for(integer i = 0; i < DEPTH; i++) begin
			mem[i] <= 0;
		end
		wr_ptr <= 0;
	end
	else begin
		en_cdr_prec <= en_cdr;	
		if(!en_cdr_prec && en_cdr && !full) begin
			mem[wr_ptr[PTR_WIDTH-1:0]] <= shift_register;
			wr_ptr <= wr_ptr + 1;
		end
		else begin
			mem[wr_ptr[PTR_WIDTH-1:0]] <= mem[wr_ptr[PTR_WIDTH-1:0]];
			
		end
	end
end

/////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////// END WRITE LOGIC ////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////


/////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////// BEGIN READ LOGIC //////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////

assign rd_en = psel && penable && !pwrite && !empty;

always_ff @(posedge clk) begin
	if(rd_en)
		prdata <= mem[rd_ptr[PTR_WIDTH-1:0]];
	else
		prdata <= 'h0;
end	

always_ff @(posedge clk, negedge reset_n) begin
	if(~reset_n) begin
		rd_ptr <= 'h0;
	end
	else begin
		if (rd_en) 
			rd_ptr <= rd_ptr + 1;
		else
			rd_ptr <= rd_ptr;
	end
end
////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////// END READ LOGIC ///////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////


endmodule



