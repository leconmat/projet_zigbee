
module zigbee_platform ( clk_i, resetn_i, mux_i, mux_o, sel_i );
  input [21:0] mux_i;
  output [17:0] mux_o;
  input [1:0] sel_i;
  input clk_i, resetn_i;
  wire   \*Logic1* , fifo_tx_pwrite_i, fifo_tx_pen_i, fifo_tx_pslv_err_o,
         fifo_tx_enable_o, fifo_tx_mem_state_o, mod_iq_enable_i, mod_iq_data_i,
         mod_iq_valid_o, demod_iq_valid_o, cordic_valid_i, cordic_valid_o,
         cdr_valid_i, cdr_valid_o, fifo_rx_valid_i, fifo_rx_data_i,
         fifo_rx_psel_i, fifo_rx_pslv_err_o, N10, N11, N12, N13, n3, n4, n5,
         n6, n7, n8, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n25, n27, n28, n29, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n73, n80, n81, \i_fifo_tx/n529 , \i_fifo_tx/n528 ,
         \i_fifo_tx/n527 , \i_fifo_tx/n526 , \i_fifo_tx/n525 ,
         \i_fifo_tx/n524 , \i_fifo_tx/n523 , \i_fifo_tx/n522 ,
         \i_fifo_tx/n521 , \i_fifo_tx/n520 , \i_fifo_tx/n519 ,
         \i_fifo_tx/n518 , \i_fifo_tx/n517 , \i_fifo_tx/n516 ,
         \i_fifo_tx/n515 , \i_fifo_tx/n514 , \i_fifo_tx/n513 ,
         \i_fifo_tx/n512 , \i_fifo_tx/n511 , \i_fifo_tx/n510 ,
         \i_fifo_tx/n509 , \i_fifo_tx/n508 , \i_fifo_tx/n507 ,
         \i_fifo_tx/n506 , \i_fifo_tx/n505 , \i_fifo_tx/n504 ,
         \i_fifo_tx/n503 , \i_fifo_tx/n502 , \i_fifo_tx/n501 ,
         \i_fifo_tx/n500 , \i_fifo_tx/n499 , \i_fifo_tx/n498 ,
         \i_fifo_tx/n497 , \i_fifo_tx/n496 , \i_fifo_tx/n495 ,
         \i_fifo_tx/n494 , \i_fifo_tx/n493 , \i_fifo_tx/n492 ,
         \i_fifo_tx/n491 , \i_fifo_tx/n490 , \i_fifo_tx/n489 ,
         \i_fifo_tx/n488 , \i_fifo_tx/n487 , \i_fifo_tx/n486 ,
         \i_fifo_tx/n485 , \i_fifo_tx/n484 , \i_fifo_tx/n483 ,
         \i_fifo_tx/n482 , \i_fifo_tx/n481 , \i_fifo_tx/n480 ,
         \i_fifo_tx/n479 , \i_fifo_tx/n478 , \i_fifo_tx/n477 ,
         \i_fifo_tx/n476 , \i_fifo_tx/n475 , \i_fifo_tx/n474 ,
         \i_fifo_tx/n473 , \i_fifo_tx/n472 , \i_fifo_tx/n471 ,
         \i_fifo_tx/n470 , \i_fifo_tx/n469 , \i_fifo_tx/n468 ,
         \i_fifo_tx/n467 , \i_fifo_tx/n466 , \i_fifo_tx/n465 ,
         \i_fifo_tx/n464 , \i_fifo_tx/n463 , \i_fifo_tx/n462 ,
         \i_fifo_tx/n461 , \i_fifo_tx/n460 , \i_fifo_tx/n459 ,
         \i_fifo_tx/n458 , \i_fifo_tx/n457 , \i_fifo_tx/n456 ,
         \i_fifo_tx/n455 , \i_fifo_tx/n454 , \i_fifo_tx/n453 ,
         \i_fifo_tx/n452 , \i_fifo_tx/n451 , \i_fifo_tx/n450 ,
         \i_fifo_tx/n449 , \i_fifo_tx/n448 , \i_fifo_tx/n447 ,
         \i_fifo_tx/n446 , \i_fifo_tx/n445 , \i_fifo_tx/n444 ,
         \i_fifo_tx/n443 , \i_fifo_tx/n442 , \i_fifo_tx/n441 ,
         \i_fifo_tx/n440 , \i_fifo_tx/n439 , \i_fifo_tx/n438 ,
         \i_fifo_tx/n437 , \i_fifo_tx/n436 , \i_fifo_tx/n435 ,
         \i_fifo_tx/n434 , \i_fifo_tx/n433 , \i_fifo_tx/n432 ,
         \i_fifo_tx/n431 , \i_fifo_tx/n430 , \i_fifo_tx/n429 ,
         \i_fifo_tx/n428 , \i_fifo_tx/n427 , \i_fifo_tx/n426 ,
         \i_fifo_tx/n425 , \i_fifo_tx/n424 , \i_fifo_tx/n423 ,
         \i_fifo_tx/n422 , \i_fifo_tx/n421 , \i_fifo_tx/n420 ,
         \i_fifo_tx/n419 , \i_fifo_tx/n418 , \i_fifo_tx/n417 ,
         \i_fifo_tx/n416 , \i_fifo_tx/n415 , \i_fifo_tx/n414 ,
         \i_fifo_tx/n413 , \i_fifo_tx/n412 , \i_fifo_tx/n411 ,
         \i_fifo_tx/n410 , \i_fifo_tx/n409 , \i_fifo_tx/n408 ,
         \i_fifo_tx/n407 , \i_fifo_tx/n406 , \i_fifo_tx/n405 ,
         \i_fifo_tx/n404 , \i_fifo_tx/n403 , \i_fifo_tx/n402 ,
         \i_fifo_tx/n401 , \i_fifo_tx/n400 , \i_fifo_tx/n399 ,
         \i_fifo_tx/n398 , \i_fifo_tx/n397 , \i_fifo_tx/n396 ,
         \i_fifo_tx/n395 , \i_fifo_tx/n394 , \i_fifo_tx/n393 ,
         \i_fifo_tx/n392 , \i_fifo_tx/n391 , \i_fifo_tx/n390 ,
         \i_fifo_tx/n389 , \i_fifo_tx/n388 , \i_fifo_tx/n387 ,
         \i_fifo_tx/n386 , \i_fifo_tx/n385 , \i_fifo_tx/n384 ,
         \i_fifo_tx/n383 , \i_fifo_tx/n382 , \i_fifo_tx/n381 ,
         \i_fifo_tx/n380 , \i_fifo_tx/n379 , \i_fifo_tx/n378 ,
         \i_fifo_tx/n377 , \i_fifo_tx/n376 , \i_fifo_tx/n375 ,
         \i_fifo_tx/n374 , \i_fifo_tx/n373 , \i_fifo_tx/n372 ,
         \i_fifo_tx/n371 , \i_fifo_tx/n370 , \i_fifo_tx/n369 ,
         \i_fifo_tx/n368 , \i_fifo_tx/n367 , \i_fifo_tx/n366 ,
         \i_fifo_tx/n365 , \i_fifo_tx/n364 , \i_fifo_tx/n363 ,
         \i_fifo_tx/n362 , \i_fifo_tx/n361 , \i_fifo_tx/n360 ,
         \i_fifo_tx/n359 , \i_fifo_tx/n358 , \i_fifo_tx/n357 ,
         \i_fifo_tx/n356 , \i_fifo_tx/n355 , \i_fifo_tx/n354 ,
         \i_fifo_tx/n353 , \i_fifo_tx/n352 , \i_fifo_tx/n351 ,
         \i_fifo_tx/n350 , \i_fifo_tx/n349 , \i_fifo_tx/n348 ,
         \i_fifo_tx/n347 , \i_fifo_tx/n346 , \i_fifo_tx/n345 ,
         \i_fifo_tx/n344 , \i_fifo_tx/n343 , \i_fifo_tx/n342 ,
         \i_fifo_tx/n341 , \i_fifo_tx/n340 , \i_fifo_tx/n339 ,
         \i_fifo_tx/n338 , \i_fifo_tx/n337 , \i_fifo_tx/n336 ,
         \i_fifo_tx/n335 , \i_fifo_tx/n334 , \i_fifo_tx/n333 ,
         \i_fifo_tx/n332 , \i_fifo_tx/n331 , \i_fifo_tx/n330 ,
         \i_fifo_tx/n329 , \i_fifo_tx/n328 , \i_fifo_tx/n327 ,
         \i_fifo_tx/n326 , \i_fifo_tx/n325 , \i_fifo_tx/n324 ,
         \i_fifo_tx/n323 , \i_fifo_tx/n322 , \i_fifo_tx/n321 ,
         \i_fifo_tx/n320 , \i_fifo_tx/n319 , \i_fifo_tx/n318 ,
         \i_fifo_tx/n317 , \i_fifo_tx/n316 , \i_fifo_tx/n315 ,
         \i_fifo_tx/n314 , \i_fifo_tx/n313 , \i_fifo_tx/n312 ,
         \i_fifo_tx/n311 , \i_fifo_tx/n310 , \i_fifo_tx/n309 ,
         \i_fifo_tx/n308 , \i_fifo_tx/n307 , \i_fifo_tx/n306 ,
         \i_fifo_tx/n305 , \i_fifo_tx/n304 , \i_fifo_tx/n303 ,
         \i_fifo_tx/n302 , \i_fifo_tx/n301 , \i_fifo_tx/n300 ,
         \i_fifo_tx/n299 , \i_fifo_tx/n298 , \i_fifo_tx/n297 ,
         \i_fifo_tx/n296 , \i_fifo_tx/n295 , \i_fifo_tx/n294 ,
         \i_fifo_tx/n293 , \i_fifo_tx/n292 , \i_fifo_tx/n291 ,
         \i_fifo_tx/n290 , \i_fifo_tx/n289 , \i_fifo_tx/n288 ,
         \i_fifo_tx/n287 , \i_fifo_tx/n286 , \i_fifo_tx/n285 ,
         \i_fifo_tx/n284 , \i_fifo_tx/n283 , \i_fifo_tx/n282 ,
         \i_fifo_tx/n281 , \i_fifo_tx/n280 , \i_fifo_tx/n279 ,
         \i_fifo_tx/n278 , \i_fifo_tx/n277 , \i_fifo_tx/n276 ,
         \i_fifo_tx/n275 , \i_fifo_tx/n274 , \i_fifo_tx/n273 ,
         \i_fifo_tx/n272 , \i_fifo_tx/n271 , \i_fifo_tx/n270 ,
         \i_fifo_tx/n269 , \i_fifo_tx/n268 , \i_fifo_tx/n267 ,
         \i_fifo_tx/n266 , \i_fifo_tx/n265 , \i_fifo_tx/n264 ,
         \i_fifo_tx/n263 , \i_fifo_tx/n262 , \i_fifo_tx/n261 ,
         \i_fifo_tx/n260 , \i_fifo_tx/n259 , \i_fifo_tx/n258 ,
         \i_fifo_tx/n257 , \i_fifo_tx/n256 , \i_fifo_tx/n255 ,
         \i_fifo_tx/n254 , \i_fifo_tx/n253 , \i_fifo_tx/n252 ,
         \i_fifo_tx/n251 , \i_fifo_tx/n250 , \i_fifo_tx/n249 ,
         \i_fifo_tx/n248 , \i_fifo_tx/n247 , \i_fifo_tx/n246 ,
         \i_fifo_tx/n245 , \i_fifo_tx/n244 , \i_fifo_tx/n243 ,
         \i_fifo_tx/n242 , \i_fifo_tx/n241 , \i_fifo_tx/n240 ,
         \i_fifo_tx/n239 , \i_fifo_tx/n238 , \i_fifo_tx/n237 ,
         \i_fifo_tx/n236 , \i_fifo_tx/n235 , \i_fifo_tx/n234 ,
         \i_fifo_tx/n233 , \i_fifo_tx/n232 , \i_fifo_tx/n231 ,
         \i_fifo_tx/n230 , \i_fifo_tx/n229 , \i_fifo_tx/n228 ,
         \i_fifo_tx/n227 , \i_fifo_tx/n226 , \i_fifo_tx/n225 ,
         \i_fifo_tx/n224 , \i_fifo_tx/n223 , \i_fifo_tx/n222 ,
         \i_fifo_tx/n221 , \i_fifo_tx/n220 , \i_fifo_tx/n219 ,
         \i_fifo_tx/n218 , \i_fifo_tx/n217 , \i_fifo_tx/n216 ,
         \i_fifo_tx/n215 , \i_fifo_tx/n214 , \i_fifo_tx/n213 ,
         \i_fifo_tx/n212 , \i_fifo_tx/n211 , \i_fifo_tx/n210 ,
         \i_fifo_tx/n209 , \i_fifo_tx/n208 , \i_fifo_tx/n207 ,
         \i_fifo_tx/n206 , \i_fifo_tx/n205 , \i_fifo_tx/n204 ,
         \i_fifo_tx/n203 , \i_fifo_tx/n201 , \i_fifo_tx/n200 ,
         \i_fifo_tx/n199 , \i_fifo_tx/n196 , \i_fifo_tx/n195 ,
         \i_fifo_tx/n194 , \i_fifo_tx/n193 , \i_fifo_tx/n192 ,
         \i_fifo_tx/n191 , \i_fifo_tx/n190 , \i_fifo_tx/n189 ,
         \i_fifo_tx/n188 , \i_fifo_tx/n187 , \i_fifo_tx/n186 ,
         \i_fifo_tx/n185 , \i_fifo_tx/n184 , \i_fifo_tx/n183 ,
         \i_fifo_tx/n182 , \i_fifo_tx/n181 , \i_fifo_tx/n180 ,
         \i_fifo_tx/n179 , \i_fifo_tx/n178 , \i_fifo_tx/n177 ,
         \i_fifo_tx/n176 , \i_fifo_tx/n175 , \i_fifo_tx/n174 ,
         \i_fifo_tx/n173 , \i_fifo_tx/n172 , \i_fifo_tx/n171 ,
         \i_fifo_tx/n170 , \i_fifo_tx/n169 , \i_fifo_tx/n168 ,
         \i_fifo_tx/n167 , \i_fifo_tx/n166 , \i_fifo_tx/n165 ,
         \i_fifo_tx/n164 , \i_fifo_tx/n163 , \i_fifo_tx/n162 ,
         \i_fifo_tx/n161 , \i_fifo_tx/n153 , \i_fifo_tx/n152 ,
         \i_fifo_tx/n151 , \i_fifo_tx/n150 , \i_fifo_tx/n149 ,
         \i_fifo_tx/n148 , \i_fifo_tx/n147 , \i_fifo_tx/n146 ,
         \i_fifo_tx/n145 , \i_fifo_tx/n144 , \i_fifo_tx/n143 ,
         \i_fifo_tx/n142 , \i_fifo_tx/n141 , \i_fifo_tx/n140 ,
         \i_fifo_tx/n139 , \i_fifo_tx/n138 , \i_fifo_tx/n137 ,
         \i_fifo_tx/n136 , \i_fifo_tx/n135 , \i_fifo_tx/n134 ,
         \i_fifo_tx/n133 , \i_fifo_tx/n132 , \i_fifo_tx/n131 ,
         \i_fifo_tx/n130 , \i_fifo_tx/n129 , \i_fifo_tx/n128 ,
         \i_fifo_tx/n127 , \i_fifo_tx/n126 , \i_fifo_tx/n125 ,
         \i_fifo_tx/n124 , \i_fifo_tx/n123 , \i_fifo_tx/n122 ,
         \i_fifo_tx/n121 , \i_fifo_tx/n120 , \i_fifo_tx/n119 ,
         \i_fifo_tx/n118 , \i_fifo_tx/n117 , \i_fifo_tx/n116 ,
         \i_fifo_tx/n115 , \i_fifo_tx/n114 , \i_fifo_tx/n113 ,
         \i_fifo_tx/n112 , \i_fifo_tx/n111 , \i_fifo_tx/n110 ,
         \i_fifo_tx/n109 , \i_fifo_tx/n108 , \i_fifo_tx/n107 ,
         \i_fifo_tx/n106 , \i_fifo_tx/n105 , \i_fifo_tx/n104 ,
         \i_fifo_tx/n103 , \i_fifo_tx/n102 , \i_fifo_tx/n101 ,
         \i_fifo_tx/n100 , \i_fifo_tx/n99 , \i_fifo_tx/n98 , \i_fifo_tx/n97 ,
         \i_fifo_tx/n96 , \i_fifo_tx/n95 , \i_fifo_tx/n94 , \i_fifo_tx/n93 ,
         \i_fifo_tx/n92 , \i_fifo_tx/n91 , \i_fifo_tx/n90 , \i_fifo_tx/n89 ,
         \i_fifo_tx/n88 , \i_fifo_tx/n86 , \i_fifo_tx/n85 , \i_fifo_tx/n84 ,
         \i_fifo_tx/n83 , \i_fifo_tx/n82 , \i_fifo_tx/n81 , \i_fifo_tx/n80 ,
         \i_fifo_tx/n79 , \i_fifo_tx/n78 , \i_fifo_tx/n74 , \i_fifo_tx/n73 ,
         \i_fifo_tx/n72 , \i_fifo_tx/n71 , \i_fifo_tx/n70 , \i_fifo_tx/n69 ,
         \i_fifo_tx/n68 , \i_fifo_tx/n67 , \i_fifo_tx/n66 , \i_fifo_tx/n65 ,
         \i_fifo_tx/n64 , \i_fifo_tx/n63 , \i_fifo_tx/n62 , \i_fifo_tx/n61 ,
         \i_fifo_tx/n60 , \i_fifo_tx/n59 , \i_fifo_tx/n58 , \i_fifo_tx/n57 ,
         \i_fifo_tx/n56 , \i_fifo_tx/n55 , \i_fifo_tx/n54 , \i_fifo_tx/n53 ,
         \i_fifo_tx/n52 , \i_fifo_tx/n51 , \i_fifo_tx/n50 , \i_fifo_tx/n49 ,
         \i_fifo_tx/n48 , \i_fifo_tx/n47 , \i_fifo_tx/n46 , \i_fifo_tx/n45 ,
         \i_fifo_tx/n44 , \i_fifo_tx/n43 , \i_fifo_tx/n42 , \i_fifo_tx/n41 ,
         \i_fifo_tx/n40 , \i_fifo_tx/n39 , \i_fifo_tx/n38 , \i_fifo_tx/n37 ,
         \i_fifo_tx/n36 , \i_fifo_tx/n35 , \i_fifo_tx/n34 , \i_fifo_tx/n33 ,
         \i_fifo_tx/n32 , \i_fifo_tx/n31 , \i_fifo_tx/n30 , \i_fifo_tx/n29 ,
         \i_fifo_tx/n28 , \i_fifo_tx/n27 , \i_fifo_tx/n26 , \i_fifo_tx/n25 ,
         \i_fifo_tx/n24 , \i_fifo_tx/n23 , \i_fifo_tx/n22 , \i_fifo_tx/n21 ,
         \i_fifo_tx/n20 , \i_fifo_tx/n19 , \i_fifo_tx/n18 , \i_fifo_tx/n17 ,
         \i_fifo_tx/n16 , \i_fifo_tx/n15 , \i_fifo_tx/n14 , \i_fifo_tx/n13 ,
         \i_fifo_tx/n12 , \i_fifo_tx/n11 , \i_fifo_tx/n10 , \i_fifo_tx/n9 ,
         \i_fifo_tx/n8 , \i_fifo_tx/n7 , \i_fifo_tx/n6 , \i_fifo_tx/n5 ,
         \i_fifo_tx/n4 , \i_fifo_tx/n3 , \i_fifo_tx/N191 , \i_fifo_tx/N190 ,
         \i_fifo_tx/N189 , \i_fifo_tx/N188 , \i_fifo_tx/N187 ,
         \i_fifo_tx/N161 , \i_fifo_tx/N160 , \i_fifo_tx/N159 ,
         \i_fifo_tx/N158 , \i_fifo_tx/N157 , \i_fifo_tx/N156 ,
         \i_fifo_tx/N151 , \i_fifo_tx/N150 , \i_fifo_tx/N149 ,
         \i_fifo_tx/N144 , \i_fifo_tx/N143 , \i_fifo_tx/N142 ,
         \i_fifo_tx/N141 , \i_fifo_tx/N140 , \i_fifo_tx/N139 ,
         \i_fifo_tx/N138 , \i_fifo_tx/N137 , \i_fifo_tx/N136 ,
         \i_fifo_tx/next_state_rd , \i_fifo_tx/state_rd , \i_fifo_tx/N134 ,
         \i_fifo_tx/N133 , \i_fifo_tx/N132 , \i_fifo_tx/N131 ,
         \i_fifo_tx/N130 , \i_fifo_tx/N129 , \i_fifo_tx/mem[63][7] ,
         \i_fifo_tx/mem[63][6] , \i_fifo_tx/mem[63][5] ,
         \i_fifo_tx/mem[63][4] , \i_fifo_tx/mem[63][3] ,
         \i_fifo_tx/mem[63][2] , \i_fifo_tx/mem[63][1] ,
         \i_fifo_tx/mem[63][0] , \i_fifo_tx/mem[62][7] ,
         \i_fifo_tx/mem[62][6] , \i_fifo_tx/mem[62][5] ,
         \i_fifo_tx/mem[62][4] , \i_fifo_tx/mem[62][3] ,
         \i_fifo_tx/mem[62][2] , \i_fifo_tx/mem[62][1] ,
         \i_fifo_tx/mem[62][0] , \i_fifo_tx/mem[61][7] ,
         \i_fifo_tx/mem[61][6] , \i_fifo_tx/mem[61][5] ,
         \i_fifo_tx/mem[61][4] , \i_fifo_tx/mem[61][3] ,
         \i_fifo_tx/mem[61][2] , \i_fifo_tx/mem[61][1] ,
         \i_fifo_tx/mem[61][0] , \i_fifo_tx/mem[60][7] ,
         \i_fifo_tx/mem[60][6] , \i_fifo_tx/mem[60][5] ,
         \i_fifo_tx/mem[60][4] , \i_fifo_tx/mem[60][3] ,
         \i_fifo_tx/mem[60][2] , \i_fifo_tx/mem[60][1] ,
         \i_fifo_tx/mem[60][0] , \i_fifo_tx/mem[59][7] ,
         \i_fifo_tx/mem[59][6] , \i_fifo_tx/mem[59][5] ,
         \i_fifo_tx/mem[59][4] , \i_fifo_tx/mem[59][3] ,
         \i_fifo_tx/mem[59][2] , \i_fifo_tx/mem[59][1] ,
         \i_fifo_tx/mem[59][0] , \i_fifo_tx/mem[58][7] ,
         \i_fifo_tx/mem[58][6] , \i_fifo_tx/mem[58][5] ,
         \i_fifo_tx/mem[58][4] , \i_fifo_tx/mem[58][3] ,
         \i_fifo_tx/mem[58][2] , \i_fifo_tx/mem[58][1] ,
         \i_fifo_tx/mem[58][0] , \i_fifo_tx/mem[57][7] ,
         \i_fifo_tx/mem[57][6] , \i_fifo_tx/mem[57][5] ,
         \i_fifo_tx/mem[57][4] , \i_fifo_tx/mem[57][3] ,
         \i_fifo_tx/mem[57][2] , \i_fifo_tx/mem[57][1] ,
         \i_fifo_tx/mem[57][0] , \i_fifo_tx/mem[56][7] ,
         \i_fifo_tx/mem[56][6] , \i_fifo_tx/mem[56][5] ,
         \i_fifo_tx/mem[56][4] , \i_fifo_tx/mem[56][3] ,
         \i_fifo_tx/mem[56][2] , \i_fifo_tx/mem[56][1] ,
         \i_fifo_tx/mem[56][0] , \i_fifo_tx/mem[55][7] ,
         \i_fifo_tx/mem[55][6] , \i_fifo_tx/mem[55][5] ,
         \i_fifo_tx/mem[55][4] , \i_fifo_tx/mem[55][3] ,
         \i_fifo_tx/mem[55][2] , \i_fifo_tx/mem[55][1] ,
         \i_fifo_tx/mem[55][0] , \i_fifo_tx/mem[54][7] ,
         \i_fifo_tx/mem[54][6] , \i_fifo_tx/mem[54][5] ,
         \i_fifo_tx/mem[54][4] , \i_fifo_tx/mem[54][3] ,
         \i_fifo_tx/mem[54][2] , \i_fifo_tx/mem[54][1] ,
         \i_fifo_tx/mem[54][0] , \i_fifo_tx/mem[53][7] ,
         \i_fifo_tx/mem[53][6] , \i_fifo_tx/mem[53][5] ,
         \i_fifo_tx/mem[53][4] , \i_fifo_tx/mem[53][3] ,
         \i_fifo_tx/mem[53][2] , \i_fifo_tx/mem[53][1] ,
         \i_fifo_tx/mem[53][0] , \i_fifo_tx/mem[52][7] ,
         \i_fifo_tx/mem[52][6] , \i_fifo_tx/mem[52][5] ,
         \i_fifo_tx/mem[52][4] , \i_fifo_tx/mem[52][3] ,
         \i_fifo_tx/mem[52][2] , \i_fifo_tx/mem[52][1] ,
         \i_fifo_tx/mem[52][0] , \i_fifo_tx/mem[51][7] ,
         \i_fifo_tx/mem[51][6] , \i_fifo_tx/mem[51][5] ,
         \i_fifo_tx/mem[51][4] , \i_fifo_tx/mem[51][3] ,
         \i_fifo_tx/mem[51][2] , \i_fifo_tx/mem[51][1] ,
         \i_fifo_tx/mem[51][0] , \i_fifo_tx/mem[50][7] ,
         \i_fifo_tx/mem[50][6] , \i_fifo_tx/mem[50][5] ,
         \i_fifo_tx/mem[50][4] , \i_fifo_tx/mem[50][3] ,
         \i_fifo_tx/mem[50][2] , \i_fifo_tx/mem[50][1] ,
         \i_fifo_tx/mem[50][0] , \i_fifo_tx/mem[49][7] ,
         \i_fifo_tx/mem[49][6] , \i_fifo_tx/mem[49][5] ,
         \i_fifo_tx/mem[49][4] , \i_fifo_tx/mem[49][3] ,
         \i_fifo_tx/mem[49][2] , \i_fifo_tx/mem[49][1] ,
         \i_fifo_tx/mem[49][0] , \i_fifo_tx/mem[48][7] ,
         \i_fifo_tx/mem[48][6] , \i_fifo_tx/mem[48][5] ,
         \i_fifo_tx/mem[48][4] , \i_fifo_tx/mem[48][3] ,
         \i_fifo_tx/mem[48][2] , \i_fifo_tx/mem[48][1] ,
         \i_fifo_tx/mem[48][0] , \i_fifo_tx/mem[47][7] ,
         \i_fifo_tx/mem[47][6] , \i_fifo_tx/mem[47][5] ,
         \i_fifo_tx/mem[47][4] , \i_fifo_tx/mem[47][3] ,
         \i_fifo_tx/mem[47][2] , \i_fifo_tx/mem[47][1] ,
         \i_fifo_tx/mem[47][0] , \i_fifo_tx/mem[46][7] ,
         \i_fifo_tx/mem[46][6] , \i_fifo_tx/mem[46][5] ,
         \i_fifo_tx/mem[46][4] , \i_fifo_tx/mem[46][3] ,
         \i_fifo_tx/mem[46][2] , \i_fifo_tx/mem[46][1] ,
         \i_fifo_tx/mem[46][0] , \i_fifo_tx/mem[45][7] ,
         \i_fifo_tx/mem[45][6] , \i_fifo_tx/mem[45][5] ,
         \i_fifo_tx/mem[45][4] , \i_fifo_tx/mem[45][3] ,
         \i_fifo_tx/mem[45][2] , \i_fifo_tx/mem[45][1] ,
         \i_fifo_tx/mem[45][0] , \i_fifo_tx/mem[44][7] ,
         \i_fifo_tx/mem[44][6] , \i_fifo_tx/mem[44][5] ,
         \i_fifo_tx/mem[44][4] , \i_fifo_tx/mem[44][3] ,
         \i_fifo_tx/mem[44][2] , \i_fifo_tx/mem[44][1] ,
         \i_fifo_tx/mem[44][0] , \i_fifo_tx/mem[43][7] ,
         \i_fifo_tx/mem[43][6] , \i_fifo_tx/mem[43][5] ,
         \i_fifo_tx/mem[43][4] , \i_fifo_tx/mem[43][3] ,
         \i_fifo_tx/mem[43][2] , \i_fifo_tx/mem[43][1] ,
         \i_fifo_tx/mem[43][0] , \i_fifo_tx/mem[42][7] ,
         \i_fifo_tx/mem[42][6] , \i_fifo_tx/mem[42][5] ,
         \i_fifo_tx/mem[42][4] , \i_fifo_tx/mem[42][3] ,
         \i_fifo_tx/mem[42][2] , \i_fifo_tx/mem[42][1] ,
         \i_fifo_tx/mem[42][0] , \i_fifo_tx/mem[41][7] ,
         \i_fifo_tx/mem[41][6] , \i_fifo_tx/mem[41][5] ,
         \i_fifo_tx/mem[41][4] , \i_fifo_tx/mem[41][3] ,
         \i_fifo_tx/mem[41][2] , \i_fifo_tx/mem[41][1] ,
         \i_fifo_tx/mem[41][0] , \i_fifo_tx/mem[40][7] ,
         \i_fifo_tx/mem[40][6] , \i_fifo_tx/mem[40][5] ,
         \i_fifo_tx/mem[40][4] , \i_fifo_tx/mem[40][3] ,
         \i_fifo_tx/mem[40][2] , \i_fifo_tx/mem[40][1] ,
         \i_fifo_tx/mem[40][0] , \i_fifo_tx/mem[39][7] ,
         \i_fifo_tx/mem[39][6] , \i_fifo_tx/mem[39][5] ,
         \i_fifo_tx/mem[39][4] , \i_fifo_tx/mem[39][3] ,
         \i_fifo_tx/mem[39][2] , \i_fifo_tx/mem[39][1] ,
         \i_fifo_tx/mem[39][0] , \i_fifo_tx/mem[38][7] ,
         \i_fifo_tx/mem[38][6] , \i_fifo_tx/mem[38][5] ,
         \i_fifo_tx/mem[38][4] , \i_fifo_tx/mem[38][3] ,
         \i_fifo_tx/mem[38][2] , \i_fifo_tx/mem[38][1] ,
         \i_fifo_tx/mem[38][0] , \i_fifo_tx/mem[37][7] ,
         \i_fifo_tx/mem[37][6] , \i_fifo_tx/mem[37][5] ,
         \i_fifo_tx/mem[37][4] , \i_fifo_tx/mem[37][3] ,
         \i_fifo_tx/mem[37][2] , \i_fifo_tx/mem[37][1] ,
         \i_fifo_tx/mem[37][0] , \i_fifo_tx/mem[36][7] ,
         \i_fifo_tx/mem[36][6] , \i_fifo_tx/mem[36][5] ,
         \i_fifo_tx/mem[36][4] , \i_fifo_tx/mem[36][3] ,
         \i_fifo_tx/mem[36][2] , \i_fifo_tx/mem[36][1] ,
         \i_fifo_tx/mem[36][0] , \i_fifo_tx/mem[35][7] ,
         \i_fifo_tx/mem[35][6] , \i_fifo_tx/mem[35][5] ,
         \i_fifo_tx/mem[35][4] , \i_fifo_tx/mem[35][3] ,
         \i_fifo_tx/mem[35][2] , \i_fifo_tx/mem[35][1] ,
         \i_fifo_tx/mem[35][0] , \i_fifo_tx/mem[34][7] ,
         \i_fifo_tx/mem[34][6] , \i_fifo_tx/mem[34][5] ,
         \i_fifo_tx/mem[34][4] , \i_fifo_tx/mem[34][3] ,
         \i_fifo_tx/mem[34][2] , \i_fifo_tx/mem[34][1] ,
         \i_fifo_tx/mem[34][0] , \i_fifo_tx/mem[33][7] ,
         \i_fifo_tx/mem[33][6] , \i_fifo_tx/mem[33][5] ,
         \i_fifo_tx/mem[33][4] , \i_fifo_tx/mem[33][3] ,
         \i_fifo_tx/mem[33][2] , \i_fifo_tx/mem[33][1] ,
         \i_fifo_tx/mem[33][0] , \i_fifo_tx/mem[32][7] ,
         \i_fifo_tx/mem[32][6] , \i_fifo_tx/mem[32][5] ,
         \i_fifo_tx/mem[32][4] , \i_fifo_tx/mem[32][3] ,
         \i_fifo_tx/mem[32][2] , \i_fifo_tx/mem[32][1] ,
         \i_fifo_tx/mem[32][0] , \i_fifo_tx/mem[31][7] ,
         \i_fifo_tx/mem[31][6] , \i_fifo_tx/mem[31][5] ,
         \i_fifo_tx/mem[31][4] , \i_fifo_tx/mem[31][3] ,
         \i_fifo_tx/mem[31][2] , \i_fifo_tx/mem[31][1] ,
         \i_fifo_tx/mem[31][0] , \i_fifo_tx/mem[30][7] ,
         \i_fifo_tx/mem[30][6] , \i_fifo_tx/mem[30][5] ,
         \i_fifo_tx/mem[30][4] , \i_fifo_tx/mem[30][3] ,
         \i_fifo_tx/mem[30][2] , \i_fifo_tx/mem[30][1] ,
         \i_fifo_tx/mem[30][0] , \i_fifo_tx/mem[29][7] ,
         \i_fifo_tx/mem[29][6] , \i_fifo_tx/mem[29][5] ,
         \i_fifo_tx/mem[29][4] , \i_fifo_tx/mem[29][3] ,
         \i_fifo_tx/mem[29][2] , \i_fifo_tx/mem[29][1] ,
         \i_fifo_tx/mem[29][0] , \i_fifo_tx/mem[28][7] ,
         \i_fifo_tx/mem[28][6] , \i_fifo_tx/mem[28][5] ,
         \i_fifo_tx/mem[28][4] , \i_fifo_tx/mem[28][3] ,
         \i_fifo_tx/mem[28][2] , \i_fifo_tx/mem[28][1] ,
         \i_fifo_tx/mem[28][0] , \i_fifo_tx/mem[27][7] ,
         \i_fifo_tx/mem[27][6] , \i_fifo_tx/mem[27][5] ,
         \i_fifo_tx/mem[27][4] , \i_fifo_tx/mem[27][3] ,
         \i_fifo_tx/mem[27][2] , \i_fifo_tx/mem[27][1] ,
         \i_fifo_tx/mem[27][0] , \i_fifo_tx/mem[26][7] ,
         \i_fifo_tx/mem[26][6] , \i_fifo_tx/mem[26][5] ,
         \i_fifo_tx/mem[26][4] , \i_fifo_tx/mem[26][3] ,
         \i_fifo_tx/mem[26][2] , \i_fifo_tx/mem[26][1] ,
         \i_fifo_tx/mem[26][0] , \i_fifo_tx/mem[25][7] ,
         \i_fifo_tx/mem[25][6] , \i_fifo_tx/mem[25][5] ,
         \i_fifo_tx/mem[25][4] , \i_fifo_tx/mem[25][3] ,
         \i_fifo_tx/mem[25][2] , \i_fifo_tx/mem[25][1] ,
         \i_fifo_tx/mem[25][0] , \i_fifo_tx/mem[24][7] ,
         \i_fifo_tx/mem[24][6] , \i_fifo_tx/mem[24][5] ,
         \i_fifo_tx/mem[24][4] , \i_fifo_tx/mem[24][3] ,
         \i_fifo_tx/mem[24][2] , \i_fifo_tx/mem[24][1] ,
         \i_fifo_tx/mem[24][0] , \i_fifo_tx/mem[23][7] ,
         \i_fifo_tx/mem[23][6] , \i_fifo_tx/mem[23][5] ,
         \i_fifo_tx/mem[23][4] , \i_fifo_tx/mem[23][3] ,
         \i_fifo_tx/mem[23][2] , \i_fifo_tx/mem[23][1] ,
         \i_fifo_tx/mem[23][0] , \i_fifo_tx/mem[22][7] ,
         \i_fifo_tx/mem[22][6] , \i_fifo_tx/mem[22][5] ,
         \i_fifo_tx/mem[22][4] , \i_fifo_tx/mem[22][3] ,
         \i_fifo_tx/mem[22][2] , \i_fifo_tx/mem[22][1] ,
         \i_fifo_tx/mem[22][0] , \i_fifo_tx/mem[21][7] ,
         \i_fifo_tx/mem[21][6] , \i_fifo_tx/mem[21][5] ,
         \i_fifo_tx/mem[21][4] , \i_fifo_tx/mem[21][3] ,
         \i_fifo_tx/mem[21][2] , \i_fifo_tx/mem[21][1] ,
         \i_fifo_tx/mem[21][0] , \i_fifo_tx/mem[20][7] ,
         \i_fifo_tx/mem[20][6] , \i_fifo_tx/mem[20][5] ,
         \i_fifo_tx/mem[20][4] , \i_fifo_tx/mem[20][3] ,
         \i_fifo_tx/mem[20][2] , \i_fifo_tx/mem[20][1] ,
         \i_fifo_tx/mem[20][0] , \i_fifo_tx/mem[19][7] ,
         \i_fifo_tx/mem[19][6] , \i_fifo_tx/mem[19][5] ,
         \i_fifo_tx/mem[19][4] , \i_fifo_tx/mem[19][3] ,
         \i_fifo_tx/mem[19][2] , \i_fifo_tx/mem[19][1] ,
         \i_fifo_tx/mem[19][0] , \i_fifo_tx/mem[18][7] ,
         \i_fifo_tx/mem[18][6] , \i_fifo_tx/mem[18][5] ,
         \i_fifo_tx/mem[18][4] , \i_fifo_tx/mem[18][3] ,
         \i_fifo_tx/mem[18][2] , \i_fifo_tx/mem[18][1] ,
         \i_fifo_tx/mem[18][0] , \i_fifo_tx/mem[17][7] ,
         \i_fifo_tx/mem[17][6] , \i_fifo_tx/mem[17][5] ,
         \i_fifo_tx/mem[17][4] , \i_fifo_tx/mem[17][3] ,
         \i_fifo_tx/mem[17][2] , \i_fifo_tx/mem[17][1] ,
         \i_fifo_tx/mem[17][0] , \i_fifo_tx/mem[16][7] ,
         \i_fifo_tx/mem[16][6] , \i_fifo_tx/mem[16][5] ,
         \i_fifo_tx/mem[16][4] , \i_fifo_tx/mem[16][3] ,
         \i_fifo_tx/mem[16][2] , \i_fifo_tx/mem[16][1] ,
         \i_fifo_tx/mem[16][0] , \i_fifo_tx/mem[15][7] ,
         \i_fifo_tx/mem[15][6] , \i_fifo_tx/mem[15][5] ,
         \i_fifo_tx/mem[15][4] , \i_fifo_tx/mem[15][3] ,
         \i_fifo_tx/mem[15][2] , \i_fifo_tx/mem[15][1] ,
         \i_fifo_tx/mem[15][0] , \i_fifo_tx/mem[14][7] ,
         \i_fifo_tx/mem[14][6] , \i_fifo_tx/mem[14][5] ,
         \i_fifo_tx/mem[14][4] , \i_fifo_tx/mem[14][3] ,
         \i_fifo_tx/mem[14][2] , \i_fifo_tx/mem[14][1] ,
         \i_fifo_tx/mem[14][0] , \i_fifo_tx/mem[13][7] ,
         \i_fifo_tx/mem[13][6] , \i_fifo_tx/mem[13][5] ,
         \i_fifo_tx/mem[13][4] , \i_fifo_tx/mem[13][3] ,
         \i_fifo_tx/mem[13][2] , \i_fifo_tx/mem[13][1] ,
         \i_fifo_tx/mem[13][0] , \i_fifo_tx/mem[12][7] ,
         \i_fifo_tx/mem[12][6] , \i_fifo_tx/mem[12][5] ,
         \i_fifo_tx/mem[12][4] , \i_fifo_tx/mem[12][3] ,
         \i_fifo_tx/mem[12][2] , \i_fifo_tx/mem[12][1] ,
         \i_fifo_tx/mem[12][0] , \i_fifo_tx/mem[11][7] ,
         \i_fifo_tx/mem[11][6] , \i_fifo_tx/mem[11][5] ,
         \i_fifo_tx/mem[11][4] , \i_fifo_tx/mem[11][3] ,
         \i_fifo_tx/mem[11][2] , \i_fifo_tx/mem[11][1] ,
         \i_fifo_tx/mem[11][0] , \i_fifo_tx/mem[10][7] ,
         \i_fifo_tx/mem[10][6] , \i_fifo_tx/mem[10][5] ,
         \i_fifo_tx/mem[10][4] , \i_fifo_tx/mem[10][3] ,
         \i_fifo_tx/mem[10][2] , \i_fifo_tx/mem[10][1] ,
         \i_fifo_tx/mem[10][0] , \i_fifo_tx/mem[9][7] , \i_fifo_tx/mem[9][6] ,
         \i_fifo_tx/mem[9][5] , \i_fifo_tx/mem[9][4] , \i_fifo_tx/mem[9][3] ,
         \i_fifo_tx/mem[9][2] , \i_fifo_tx/mem[9][1] , \i_fifo_tx/mem[9][0] ,
         \i_fifo_tx/mem[8][7] , \i_fifo_tx/mem[8][6] , \i_fifo_tx/mem[8][5] ,
         \i_fifo_tx/mem[8][4] , \i_fifo_tx/mem[8][3] , \i_fifo_tx/mem[8][2] ,
         \i_fifo_tx/mem[8][1] , \i_fifo_tx/mem[8][0] , \i_fifo_tx/mem[7][7] ,
         \i_fifo_tx/mem[7][6] , \i_fifo_tx/mem[7][5] , \i_fifo_tx/mem[7][4] ,
         \i_fifo_tx/mem[7][3] , \i_fifo_tx/mem[7][2] , \i_fifo_tx/mem[7][1] ,
         \i_fifo_tx/mem[7][0] , \i_fifo_tx/mem[6][7] , \i_fifo_tx/mem[6][6] ,
         \i_fifo_tx/mem[6][5] , \i_fifo_tx/mem[6][4] , \i_fifo_tx/mem[6][3] ,
         \i_fifo_tx/mem[6][2] , \i_fifo_tx/mem[6][1] , \i_fifo_tx/mem[6][0] ,
         \i_fifo_tx/mem[5][7] , \i_fifo_tx/mem[5][6] , \i_fifo_tx/mem[5][5] ,
         \i_fifo_tx/mem[5][4] , \i_fifo_tx/mem[5][3] , \i_fifo_tx/mem[5][2] ,
         \i_fifo_tx/mem[5][1] , \i_fifo_tx/mem[5][0] , \i_fifo_tx/mem[4][7] ,
         \i_fifo_tx/mem[4][6] , \i_fifo_tx/mem[4][5] , \i_fifo_tx/mem[4][4] ,
         \i_fifo_tx/mem[4][3] , \i_fifo_tx/mem[4][2] , \i_fifo_tx/mem[4][1] ,
         \i_fifo_tx/mem[4][0] , \i_fifo_tx/mem[3][7] , \i_fifo_tx/mem[3][6] ,
         \i_fifo_tx/mem[3][5] , \i_fifo_tx/mem[3][4] , \i_fifo_tx/mem[3][3] ,
         \i_fifo_tx/mem[3][2] , \i_fifo_tx/mem[3][1] , \i_fifo_tx/mem[3][0] ,
         \i_fifo_tx/mem[2][7] , \i_fifo_tx/mem[2][6] , \i_fifo_tx/mem[2][5] ,
         \i_fifo_tx/mem[2][4] , \i_fifo_tx/mem[2][3] , \i_fifo_tx/mem[2][2] ,
         \i_fifo_tx/mem[2][1] , \i_fifo_tx/mem[2][0] , \i_fifo_tx/mem[1][7] ,
         \i_fifo_tx/mem[1][6] , \i_fifo_tx/mem[1][5] , \i_fifo_tx/mem[1][4] ,
         \i_fifo_tx/mem[1][3] , \i_fifo_tx/mem[1][2] , \i_fifo_tx/mem[1][1] ,
         \i_fifo_tx/mem[1][0] , \i_fifo_tx/mem[0][7] , \i_fifo_tx/mem[0][6] ,
         \i_fifo_tx/mem[0][5] , \i_fifo_tx/mem[0][4] , \i_fifo_tx/mem[0][3] ,
         \i_fifo_tx/mem[0][2] , \i_fifo_tx/mem[0][1] , \i_fifo_tx/mem[0][0] ,
         \i_fifo_tx/N40 , \i_fifo_tx/rd_ptr[6] , \i_fifo_tx/wr_ptr[6] ,
         \i_fifo_tx/N38 , \i_fifo_tx/N37 , \i_fifo_tx/N36 , \i_fifo_tx/N35 ,
         \i_fifo_tx/N34 , \i_fifo_tx/N33 , \i_fifo_tx/N32 , \i_fifo_tx/N31 ,
         \i_fifo_tx/N30 , \i_fifo_tx/N29 , \i_fifo_tx/N28 , \i_fifo_tx/N27 ,
         \i_fifo_tx/N26 , \i_mod_iq/en_10MHz , \i_iq_demod/filter_en ,
         \i_cordic/n22 , \i_cordic/n21 , \i_cordic/n20 , \i_cordic/n19 ,
         \i_cordic/n16 , \i_cordic/n14 , \i_cordic/n12 , \i_cordic/n10 ,
         \i_cordic/n7 , \i_cordic/n6 , \i_cordic/n5 , \i_cordic/N16 ,
         \i_cordic/N15 , \i_cordic/N14 , \i_cordic/N13 , \i_cordic/N10 ,
         \i_cordic/N9 , \i_cordic/N8 , \i_cordic/N7 , \i_cordic/N6 ,
         \i_cordic/valid_s1[4] , \i_cordic/cor_w_s1[4][5] ,
         \i_cordic/cor_w_s1[4][4] , \i_cordic/cor_w_s1[4][3] ,
         \i_cordic/cor_w_s1[4][2] , \i_cordic/cor_y_s1[2][5] ,
         \i_cordic/cor_y_s1[2][4] , \i_cordic/cor_y_s1[2][3] ,
         \i_cordic/cor_y_s1[2][2] , \i_cordic/cor_y_s1[2][1] ,
         \i_cordic/cor_x_s1[2][5] , \i_cordic/cor_x_s1[2][4] ,
         \i_cordic/cor_x_s1[2][3] , \i_cordic/cor_x_s1[2][2] ,
         \i_cordic/valid_s0[2] , \i_cordic/cor_w_s0[2][4] ,
         \i_cordic/cor_w_s0[2][5] , \i_cordic/cor_y_s0[2][5] ,
         \i_cordic/cor_y_s0[2][4] , \i_cordic/cor_y_s0[2][3] ,
         \i_cordic/cor_y_s0[2][2] , \i_cordic/cor_y_s0[2][1] ,
         \i_cordic/cor_y_s0[2][0] , \i_cordic/cor_y_s0[1][5] ,
         \i_cordic/cor_y_s0[1][4] , \i_cordic/cor_y_s0[1][3] ,
         \i_cordic/cor_y_s0[1][2] , \i_cordic/cor_y_s0[1][1] ,
         \i_cordic/cor_y_s0[1][0] , \i_cordic/cor_y_s0[0][5] ,
         \i_cordic/cor_y_s0[0][4] , \i_cordic/cor_y_s0[0][3] ,
         \i_cordic/cor_y_s0[0][2] , \i_cordic/cor_y_s0[0][1] ,
         \i_cordic/cor_y_s0[0][0] , \i_cordic/cor_x_s0[0][0] ,
         \i_cordic/cor_x_s0[0][1] , \i_cordic/cor_x_s0[0][2] ,
         \i_cordic/cor_x_s0[0][3] , \i_cordic/cor_x_s0[1][0] ,
         \i_cordic/cor_x_s0[1][1] , \i_cordic/cor_x_s0[1][2] ,
         \i_cordic/cor_x_s0[1][3] , \i_cordic/cor_x_s0[1][4] ,
         \i_cordic/cor_x_s0[1][5] , \i_cordic/cor_x_s0[2][2] ,
         \i_cordic/cor_x_s0[2][3] , \i_cordic/cor_x_s0[2][4] ,
         \i_cordic/cor_x_s0[2][5] , \i_cdr/data_w , \i_fifo_rx/n537 ,
         \i_fifo_rx/n536 , \i_fifo_rx/n535 , \i_fifo_rx/n534 ,
         \i_fifo_rx/n533 , \i_fifo_rx/n532 , \i_fifo_rx/n531 ,
         \i_fifo_rx/n530 , \i_fifo_rx/n529 , \i_fifo_rx/n528 ,
         \i_fifo_rx/n527 , \i_fifo_rx/n526 , \i_fifo_rx/n525 ,
         \i_fifo_rx/n524 , \i_fifo_rx/n523 , \i_fifo_rx/n522 ,
         \i_fifo_rx/n521 , \i_fifo_rx/n520 , \i_fifo_rx/n519 ,
         \i_fifo_rx/n518 , \i_fifo_rx/n517 , \i_fifo_rx/n516 ,
         \i_fifo_rx/n515 , \i_fifo_rx/n514 , \i_fifo_rx/n513 ,
         \i_fifo_rx/n512 , \i_fifo_rx/n511 , \i_fifo_rx/n510 ,
         \i_fifo_rx/n509 , \i_fifo_rx/n508 , \i_fifo_rx/n507 ,
         \i_fifo_rx/n506 , \i_fifo_rx/n505 , \i_fifo_rx/n504 ,
         \i_fifo_rx/n503 , \i_fifo_rx/n502 , \i_fifo_rx/n501 ,
         \i_fifo_rx/n500 , \i_fifo_rx/n499 , \i_fifo_rx/n498 ,
         \i_fifo_rx/n497 , \i_fifo_rx/n496 , \i_fifo_rx/n495 ,
         \i_fifo_rx/n494 , \i_fifo_rx/n493 , \i_fifo_rx/n492 ,
         \i_fifo_rx/n491 , \i_fifo_rx/n490 , \i_fifo_rx/n489 ,
         \i_fifo_rx/n488 , \i_fifo_rx/n487 , \i_fifo_rx/n486 ,
         \i_fifo_rx/n485 , \i_fifo_rx/n484 , \i_fifo_rx/n483 ,
         \i_fifo_rx/n482 , \i_fifo_rx/n481 , \i_fifo_rx/n480 ,
         \i_fifo_rx/n479 , \i_fifo_rx/n478 , \i_fifo_rx/n477 ,
         \i_fifo_rx/n476 , \i_fifo_rx/n475 , \i_fifo_rx/n474 ,
         \i_fifo_rx/n473 , \i_fifo_rx/n472 , \i_fifo_rx/n471 ,
         \i_fifo_rx/n470 , \i_fifo_rx/n469 , \i_fifo_rx/n468 ,
         \i_fifo_rx/n467 , \i_fifo_rx/n466 , \i_fifo_rx/n465 ,
         \i_fifo_rx/n464 , \i_fifo_rx/n463 , \i_fifo_rx/n462 ,
         \i_fifo_rx/n461 , \i_fifo_rx/n460 , \i_fifo_rx/n459 ,
         \i_fifo_rx/n458 , \i_fifo_rx/n457 , \i_fifo_rx/n456 ,
         \i_fifo_rx/n455 , \i_fifo_rx/n454 , \i_fifo_rx/n453 ,
         \i_fifo_rx/n452 , \i_fifo_rx/n451 , \i_fifo_rx/n450 ,
         \i_fifo_rx/n449 , \i_fifo_rx/n448 , \i_fifo_rx/n447 ,
         \i_fifo_rx/n446 , \i_fifo_rx/n445 , \i_fifo_rx/n444 ,
         \i_fifo_rx/n443 , \i_fifo_rx/n442 , \i_fifo_rx/n441 ,
         \i_fifo_rx/n440 , \i_fifo_rx/n439 , \i_fifo_rx/n438 ,
         \i_fifo_rx/n437 , \i_fifo_rx/n436 , \i_fifo_rx/n435 ,
         \i_fifo_rx/n434 , \i_fifo_rx/n433 , \i_fifo_rx/n432 ,
         \i_fifo_rx/n431 , \i_fifo_rx/n430 , \i_fifo_rx/n429 ,
         \i_fifo_rx/n428 , \i_fifo_rx/n427 , \i_fifo_rx/n426 ,
         \i_fifo_rx/n425 , \i_fifo_rx/n424 , \i_fifo_rx/n423 ,
         \i_fifo_rx/n422 , \i_fifo_rx/n421 , \i_fifo_rx/n420 ,
         \i_fifo_rx/n419 , \i_fifo_rx/n418 , \i_fifo_rx/n417 ,
         \i_fifo_rx/n416 , \i_fifo_rx/n415 , \i_fifo_rx/n414 ,
         \i_fifo_rx/n413 , \i_fifo_rx/n412 , \i_fifo_rx/n411 ,
         \i_fifo_rx/n410 , \i_fifo_rx/n409 , \i_fifo_rx/n408 ,
         \i_fifo_rx/n407 , \i_fifo_rx/n406 , \i_fifo_rx/n405 ,
         \i_fifo_rx/n404 , \i_fifo_rx/n403 , \i_fifo_rx/n402 ,
         \i_fifo_rx/n401 , \i_fifo_rx/n400 , \i_fifo_rx/n399 ,
         \i_fifo_rx/n398 , \i_fifo_rx/n397 , \i_fifo_rx/n396 ,
         \i_fifo_rx/n395 , \i_fifo_rx/n394 , \i_fifo_rx/n393 ,
         \i_fifo_rx/n392 , \i_fifo_rx/n391 , \i_fifo_rx/n390 ,
         \i_fifo_rx/n389 , \i_fifo_rx/n388 , \i_fifo_rx/n387 ,
         \i_fifo_rx/n386 , \i_fifo_rx/n385 , \i_fifo_rx/n384 ,
         \i_fifo_rx/n383 , \i_fifo_rx/n382 , \i_fifo_rx/n381 ,
         \i_fifo_rx/n380 , \i_fifo_rx/n379 , \i_fifo_rx/n378 ,
         \i_fifo_rx/n377 , \i_fifo_rx/n376 , \i_fifo_rx/n375 ,
         \i_fifo_rx/n374 , \i_fifo_rx/n373 , \i_fifo_rx/n372 ,
         \i_fifo_rx/n371 , \i_fifo_rx/n370 , \i_fifo_rx/n369 ,
         \i_fifo_rx/n368 , \i_fifo_rx/n367 , \i_fifo_rx/n366 ,
         \i_fifo_rx/n365 , \i_fifo_rx/n364 , \i_fifo_rx/n363 ,
         \i_fifo_rx/n362 , \i_fifo_rx/n361 , \i_fifo_rx/n360 ,
         \i_fifo_rx/n359 , \i_fifo_rx/n358 , \i_fifo_rx/n357 ,
         \i_fifo_rx/n356 , \i_fifo_rx/n355 , \i_fifo_rx/n354 ,
         \i_fifo_rx/n353 , \i_fifo_rx/n352 , \i_fifo_rx/n351 ,
         \i_fifo_rx/n350 , \i_fifo_rx/n349 , \i_fifo_rx/n348 ,
         \i_fifo_rx/n347 , \i_fifo_rx/n346 , \i_fifo_rx/n345 ,
         \i_fifo_rx/n344 , \i_fifo_rx/n343 , \i_fifo_rx/n342 ,
         \i_fifo_rx/n341 , \i_fifo_rx/n340 , \i_fifo_rx/n339 ,
         \i_fifo_rx/n338 , \i_fifo_rx/n337 , \i_fifo_rx/n336 ,
         \i_fifo_rx/n335 , \i_fifo_rx/n334 , \i_fifo_rx/n333 ,
         \i_fifo_rx/n332 , \i_fifo_rx/n331 , \i_fifo_rx/n330 ,
         \i_fifo_rx/n329 , \i_fifo_rx/n328 , \i_fifo_rx/n327 ,
         \i_fifo_rx/n326 , \i_fifo_rx/n325 , \i_fifo_rx/n324 ,
         \i_fifo_rx/n323 , \i_fifo_rx/n322 , \i_fifo_rx/n321 ,
         \i_fifo_rx/n320 , \i_fifo_rx/n319 , \i_fifo_rx/n318 ,
         \i_fifo_rx/n317 , \i_fifo_rx/n316 , \i_fifo_rx/n315 ,
         \i_fifo_rx/n314 , \i_fifo_rx/n313 , \i_fifo_rx/n312 ,
         \i_fifo_rx/n311 , \i_fifo_rx/n310 , \i_fifo_rx/n309 ,
         \i_fifo_rx/n308 , \i_fifo_rx/n307 , \i_fifo_rx/n306 ,
         \i_fifo_rx/n305 , \i_fifo_rx/n304 , \i_fifo_rx/n303 ,
         \i_fifo_rx/n302 , \i_fifo_rx/n301 , \i_fifo_rx/n300 ,
         \i_fifo_rx/n299 , \i_fifo_rx/n298 , \i_fifo_rx/n297 ,
         \i_fifo_rx/n296 , \i_fifo_rx/n295 , \i_fifo_rx/n294 ,
         \i_fifo_rx/n293 , \i_fifo_rx/n292 , \i_fifo_rx/n291 ,
         \i_fifo_rx/n290 , \i_fifo_rx/n289 , \i_fifo_rx/n288 ,
         \i_fifo_rx/n287 , \i_fifo_rx/n286 , \i_fifo_rx/n285 ,
         \i_fifo_rx/n284 , \i_fifo_rx/n283 , \i_fifo_rx/n282 ,
         \i_fifo_rx/n281 , \i_fifo_rx/n280 , \i_fifo_rx/n279 ,
         \i_fifo_rx/n278 , \i_fifo_rx/n277 , \i_fifo_rx/n276 ,
         \i_fifo_rx/n275 , \i_fifo_rx/n274 , \i_fifo_rx/n273 ,
         \i_fifo_rx/n272 , \i_fifo_rx/n271 , \i_fifo_rx/n270 ,
         \i_fifo_rx/n269 , \i_fifo_rx/n268 , \i_fifo_rx/n267 ,
         \i_fifo_rx/n266 , \i_fifo_rx/n265 , \i_fifo_rx/n264 ,
         \i_fifo_rx/n263 , \i_fifo_rx/n262 , \i_fifo_rx/n261 ,
         \i_fifo_rx/n260 , \i_fifo_rx/n259 , \i_fifo_rx/n258 ,
         \i_fifo_rx/n257 , \i_fifo_rx/n256 , \i_fifo_rx/n255 ,
         \i_fifo_rx/n254 , \i_fifo_rx/n253 , \i_fifo_rx/n252 ,
         \i_fifo_rx/n251 , \i_fifo_rx/n250 , \i_fifo_rx/n249 ,
         \i_fifo_rx/n248 , \i_fifo_rx/n247 , \i_fifo_rx/n246 ,
         \i_fifo_rx/n245 , \i_fifo_rx/n244 , \i_fifo_rx/n243 ,
         \i_fifo_rx/n242 , \i_fifo_rx/n241 , \i_fifo_rx/n240 ,
         \i_fifo_rx/n239 , \i_fifo_rx/n238 , \i_fifo_rx/n237 ,
         \i_fifo_rx/n236 , \i_fifo_rx/n235 , \i_fifo_rx/n234 ,
         \i_fifo_rx/n233 , \i_fifo_rx/n232 , \i_fifo_rx/n231 ,
         \i_fifo_rx/n230 , \i_fifo_rx/n229 , \i_fifo_rx/n228 ,
         \i_fifo_rx/n227 , \i_fifo_rx/n226 , \i_fifo_rx/n225 ,
         \i_fifo_rx/n224 , \i_fifo_rx/n223 , \i_fifo_rx/n222 ,
         \i_fifo_rx/n221 , \i_fifo_rx/n220 , \i_fifo_rx/n219 ,
         \i_fifo_rx/n218 , \i_fifo_rx/n217 , \i_fifo_rx/n214 ,
         \i_fifo_rx/n213 , \i_fifo_rx/n212 , \i_fifo_rx/n211 ,
         \i_fifo_rx/n210 , \i_fifo_rx/n209 , \i_fifo_rx/n198 ,
         \i_fifo_rx/n196 , \i_fifo_rx/n194 , \i_fifo_rx/n192 ,
         \i_fifo_rx/n189 , \i_fifo_rx/n188 , \i_fifo_rx/n186 ,
         \i_fifo_rx/n184 , \i_fifo_rx/n182 , \i_fifo_rx/n180 ,
         \i_fifo_rx/n179 , \i_fifo_rx/n177 , \i_fifo_rx/n176 ,
         \i_fifo_rx/n175 , \i_fifo_rx/n174 , \i_fifo_rx/n173 ,
         \i_fifo_rx/n172 , \i_fifo_rx/n171 , \i_fifo_rx/n170 ,
         \i_fifo_rx/n169 , \i_fifo_rx/n168 , \i_fifo_rx/n167 ,
         \i_fifo_rx/n166 , \i_fifo_rx/n165 , \i_fifo_rx/n164 ,
         \i_fifo_rx/n163 , \i_fifo_rx/n162 , \i_fifo_rx/n161 ,
         \i_fifo_rx/n160 , \i_fifo_rx/n159 , \i_fifo_rx/n158 ,
         \i_fifo_rx/n157 , \i_fifo_rx/n156 , \i_fifo_rx/n155 ,
         \i_fifo_rx/n154 , \i_fifo_rx/n153 , \i_fifo_rx/n152 ,
         \i_fifo_rx/n151 , \i_fifo_rx/n150 , \i_fifo_rx/n149 ,
         \i_fifo_rx/n148 , \i_fifo_rx/n147 , \i_fifo_rx/n146 ,
         \i_fifo_rx/n145 , \i_fifo_rx/n144 , \i_fifo_rx/n143 ,
         \i_fifo_rx/n142 , \i_fifo_rx/n141 , \i_fifo_rx/n140 ,
         \i_fifo_rx/n139 , \i_fifo_rx/n138 , \i_fifo_rx/n137 ,
         \i_fifo_rx/n136 , \i_fifo_rx/n135 , \i_fifo_rx/n134 ,
         \i_fifo_rx/n133 , \i_fifo_rx/n132 , \i_fifo_rx/n131 ,
         \i_fifo_rx/n130 , \i_fifo_rx/n129 , \i_fifo_rx/n128 ,
         \i_fifo_rx/n127 , \i_fifo_rx/n126 , \i_fifo_rx/n125 ,
         \i_fifo_rx/n124 , \i_fifo_rx/n123 , \i_fifo_rx/n122 ,
         \i_fifo_rx/n121 , \i_fifo_rx/n120 , \i_fifo_rx/n119 ,
         \i_fifo_rx/n118 , \i_fifo_rx/n117 , \i_fifo_rx/n116 ,
         \i_fifo_rx/n115 , \i_fifo_rx/n114 , \i_fifo_rx/n113 ,
         \i_fifo_rx/n112 , \i_fifo_rx/n111 , \i_fifo_rx/n110 ,
         \i_fifo_rx/n109 , \i_fifo_rx/n108 , \i_fifo_rx/n107 ,
         \i_fifo_rx/n106 , \i_fifo_rx/n105 , \i_fifo_rx/n104 ,
         \i_fifo_rx/n103 , \i_fifo_rx/n102 , \i_fifo_rx/n101 ,
         \i_fifo_rx/n100 , \i_fifo_rx/n99 , \i_fifo_rx/n98 , \i_fifo_rx/n97 ,
         \i_fifo_rx/n96 , \i_fifo_rx/n95 , \i_fifo_rx/n94 , \i_fifo_rx/n93 ,
         \i_fifo_rx/n92 , \i_fifo_rx/n91 , \i_fifo_rx/n90 , \i_fifo_rx/n89 ,
         \i_fifo_rx/n88 , \i_fifo_rx/n87 , \i_fifo_rx/n86 , \i_fifo_rx/n85 ,
         \i_fifo_rx/n84 , \i_fifo_rx/n83 , \i_fifo_rx/n82 , \i_fifo_rx/n81 ,
         \i_fifo_rx/n80 , \i_fifo_rx/n79 , \i_fifo_rx/n78 , \i_fifo_rx/n77 ,
         \i_fifo_rx/n76 , \i_fifo_rx/n75 , \i_fifo_rx/n74 , \i_fifo_rx/n73 ,
         \i_fifo_rx/n72 , \i_fifo_rx/n71 , \i_fifo_rx/n70 , \i_fifo_rx/n69 ,
         \i_fifo_rx/n68 , \i_fifo_rx/n67 , \i_fifo_rx/n66 , \i_fifo_rx/n65 ,
         \i_fifo_rx/n64 , \i_fifo_rx/n63 , \i_fifo_rx/n62 , \i_fifo_rx/n61 ,
         \i_fifo_rx/n60 , \i_fifo_rx/n59 , \i_fifo_rx/n58 , \i_fifo_rx/n57 ,
         \i_fifo_rx/n56 , \i_fifo_rx/n55 , \i_fifo_rx/n54 , \i_fifo_rx/n53 ,
         \i_fifo_rx/n52 , \i_fifo_rx/n51 , \i_fifo_rx/n50 , \i_fifo_rx/n49 ,
         \i_fifo_rx/n48 , \i_fifo_rx/n47 , \i_fifo_rx/n46 , \i_fifo_rx/n45 ,
         \i_fifo_rx/n44 , \i_fifo_rx/n43 , \i_fifo_rx/n42 , \i_fifo_rx/n41 ,
         \i_fifo_rx/n40 , \i_fifo_rx/n39 , \i_fifo_rx/n38 , \i_fifo_rx/n37 ,
         \i_fifo_rx/n36 , \i_fifo_rx/n35 , \i_fifo_rx/n34 , \i_fifo_rx/n33 ,
         \i_fifo_rx/n32 , \i_fifo_rx/n31 , \i_fifo_rx/n30 , \i_fifo_rx/n29 ,
         \i_fifo_rx/n28 , \i_fifo_rx/n27 , \i_fifo_rx/n26 , \i_fifo_rx/n25 ,
         \i_fifo_rx/n24 , \i_fifo_rx/n23 , \i_fifo_rx/n22 , \i_fifo_rx/n14 ,
         \i_fifo_rx/n12 , \i_fifo_rx/n11 , \i_fifo_rx/n10 , \i_fifo_rx/n9 ,
         \i_fifo_rx/n8 , \i_fifo_rx/n7 , \i_fifo_rx/n6 , \i_fifo_rx/n5 ,
         \i_fifo_rx/n4 , \i_fifo_rx/n3 , \i_fifo_rx/N694 , \i_fifo_rx/N693 ,
         \i_fifo_rx/N692 , \i_fifo_rx/N691 , \i_fifo_rx/N690 ,
         \i_fifo_rx/N689 , \i_fifo_rx/N687 , \i_fifo_rx/N686 ,
         \i_fifo_rx/N685 , \i_fifo_rx/N684 , \i_fifo_rx/N683 ,
         \i_fifo_rx/N682 , \i_fifo_rx/N681 , \i_fifo_rx/N680 , \i_fifo_rx/N94 ,
         \i_fifo_rx/N93 , \i_fifo_rx/N92 , \i_fifo_rx/N91 , \i_fifo_rx/N90 ,
         \i_fifo_rx/N89 , \i_fifo_rx/N88 , \i_fifo_rx/N87 , \i_fifo_rx/N86 ,
         \i_fifo_rx/N85 , \i_fifo_rx/N84 , \i_fifo_rx/N83 , \i_fifo_rx/N82 ,
         \i_fifo_rx/N81 , \i_fifo_rx/mem[63][7] , \i_fifo_rx/mem[63][6] ,
         \i_fifo_rx/mem[63][5] , \i_fifo_rx/mem[63][4] ,
         \i_fifo_rx/mem[63][3] , \i_fifo_rx/mem[63][2] ,
         \i_fifo_rx/mem[63][1] , \i_fifo_rx/mem[63][0] ,
         \i_fifo_rx/mem[62][7] , \i_fifo_rx/mem[62][6] ,
         \i_fifo_rx/mem[62][5] , \i_fifo_rx/mem[62][4] ,
         \i_fifo_rx/mem[62][3] , \i_fifo_rx/mem[62][2] ,
         \i_fifo_rx/mem[62][1] , \i_fifo_rx/mem[62][0] ,
         \i_fifo_rx/mem[61][7] , \i_fifo_rx/mem[61][6] ,
         \i_fifo_rx/mem[61][5] , \i_fifo_rx/mem[61][4] ,
         \i_fifo_rx/mem[61][3] , \i_fifo_rx/mem[61][2] ,
         \i_fifo_rx/mem[61][1] , \i_fifo_rx/mem[61][0] ,
         \i_fifo_rx/mem[60][7] , \i_fifo_rx/mem[60][6] ,
         \i_fifo_rx/mem[60][5] , \i_fifo_rx/mem[60][4] ,
         \i_fifo_rx/mem[60][3] , \i_fifo_rx/mem[60][2] ,
         \i_fifo_rx/mem[60][1] , \i_fifo_rx/mem[60][0] ,
         \i_fifo_rx/mem[59][7] , \i_fifo_rx/mem[59][6] ,
         \i_fifo_rx/mem[59][5] , \i_fifo_rx/mem[59][4] ,
         \i_fifo_rx/mem[59][3] , \i_fifo_rx/mem[59][2] ,
         \i_fifo_rx/mem[59][1] , \i_fifo_rx/mem[59][0] ,
         \i_fifo_rx/mem[58][7] , \i_fifo_rx/mem[58][6] ,
         \i_fifo_rx/mem[58][5] , \i_fifo_rx/mem[58][4] ,
         \i_fifo_rx/mem[58][3] , \i_fifo_rx/mem[58][2] ,
         \i_fifo_rx/mem[58][1] , \i_fifo_rx/mem[58][0] ,
         \i_fifo_rx/mem[57][7] , \i_fifo_rx/mem[57][6] ,
         \i_fifo_rx/mem[57][5] , \i_fifo_rx/mem[57][4] ,
         \i_fifo_rx/mem[57][3] , \i_fifo_rx/mem[57][2] ,
         \i_fifo_rx/mem[57][1] , \i_fifo_rx/mem[57][0] ,
         \i_fifo_rx/mem[56][7] , \i_fifo_rx/mem[56][6] ,
         \i_fifo_rx/mem[56][5] , \i_fifo_rx/mem[56][4] ,
         \i_fifo_rx/mem[56][3] , \i_fifo_rx/mem[56][2] ,
         \i_fifo_rx/mem[56][1] , \i_fifo_rx/mem[56][0] ,
         \i_fifo_rx/mem[55][7] , \i_fifo_rx/mem[55][6] ,
         \i_fifo_rx/mem[55][5] , \i_fifo_rx/mem[55][4] ,
         \i_fifo_rx/mem[55][3] , \i_fifo_rx/mem[55][2] ,
         \i_fifo_rx/mem[55][1] , \i_fifo_rx/mem[55][0] ,
         \i_fifo_rx/mem[54][7] , \i_fifo_rx/mem[54][6] ,
         \i_fifo_rx/mem[54][5] , \i_fifo_rx/mem[54][4] ,
         \i_fifo_rx/mem[54][3] , \i_fifo_rx/mem[54][2] ,
         \i_fifo_rx/mem[54][1] , \i_fifo_rx/mem[54][0] ,
         \i_fifo_rx/mem[53][7] , \i_fifo_rx/mem[53][6] ,
         \i_fifo_rx/mem[53][5] , \i_fifo_rx/mem[53][4] ,
         \i_fifo_rx/mem[53][3] , \i_fifo_rx/mem[53][2] ,
         \i_fifo_rx/mem[53][1] , \i_fifo_rx/mem[53][0] ,
         \i_fifo_rx/mem[52][7] , \i_fifo_rx/mem[52][6] ,
         \i_fifo_rx/mem[52][5] , \i_fifo_rx/mem[52][4] ,
         \i_fifo_rx/mem[52][3] , \i_fifo_rx/mem[52][2] ,
         \i_fifo_rx/mem[52][1] , \i_fifo_rx/mem[52][0] ,
         \i_fifo_rx/mem[51][7] , \i_fifo_rx/mem[51][6] ,
         \i_fifo_rx/mem[51][5] , \i_fifo_rx/mem[51][4] ,
         \i_fifo_rx/mem[51][3] , \i_fifo_rx/mem[51][2] ,
         \i_fifo_rx/mem[51][1] , \i_fifo_rx/mem[51][0] ,
         \i_fifo_rx/mem[50][7] , \i_fifo_rx/mem[50][6] ,
         \i_fifo_rx/mem[50][5] , \i_fifo_rx/mem[50][4] ,
         \i_fifo_rx/mem[50][3] , \i_fifo_rx/mem[50][2] ,
         \i_fifo_rx/mem[50][1] , \i_fifo_rx/mem[50][0] ,
         \i_fifo_rx/mem[49][7] , \i_fifo_rx/mem[49][6] ,
         \i_fifo_rx/mem[49][5] , \i_fifo_rx/mem[49][4] ,
         \i_fifo_rx/mem[49][3] , \i_fifo_rx/mem[49][2] ,
         \i_fifo_rx/mem[49][1] , \i_fifo_rx/mem[49][0] ,
         \i_fifo_rx/mem[48][7] , \i_fifo_rx/mem[48][6] ,
         \i_fifo_rx/mem[48][5] , \i_fifo_rx/mem[48][4] ,
         \i_fifo_rx/mem[48][3] , \i_fifo_rx/mem[48][2] ,
         \i_fifo_rx/mem[48][1] , \i_fifo_rx/mem[48][0] ,
         \i_fifo_rx/mem[47][7] , \i_fifo_rx/mem[47][6] ,
         \i_fifo_rx/mem[47][5] , \i_fifo_rx/mem[47][4] ,
         \i_fifo_rx/mem[47][3] , \i_fifo_rx/mem[47][2] ,
         \i_fifo_rx/mem[47][1] , \i_fifo_rx/mem[47][0] ,
         \i_fifo_rx/mem[46][7] , \i_fifo_rx/mem[46][6] ,
         \i_fifo_rx/mem[46][5] , \i_fifo_rx/mem[46][4] ,
         \i_fifo_rx/mem[46][3] , \i_fifo_rx/mem[46][2] ,
         \i_fifo_rx/mem[46][1] , \i_fifo_rx/mem[46][0] ,
         \i_fifo_rx/mem[45][7] , \i_fifo_rx/mem[45][6] ,
         \i_fifo_rx/mem[45][5] , \i_fifo_rx/mem[45][4] ,
         \i_fifo_rx/mem[45][3] , \i_fifo_rx/mem[45][2] ,
         \i_fifo_rx/mem[45][1] , \i_fifo_rx/mem[45][0] ,
         \i_fifo_rx/mem[44][7] , \i_fifo_rx/mem[44][6] ,
         \i_fifo_rx/mem[44][5] , \i_fifo_rx/mem[44][4] ,
         \i_fifo_rx/mem[44][3] , \i_fifo_rx/mem[44][2] ,
         \i_fifo_rx/mem[44][1] , \i_fifo_rx/mem[44][0] ,
         \i_fifo_rx/mem[43][7] , \i_fifo_rx/mem[43][6] ,
         \i_fifo_rx/mem[43][5] , \i_fifo_rx/mem[43][4] ,
         \i_fifo_rx/mem[43][3] , \i_fifo_rx/mem[43][2] ,
         \i_fifo_rx/mem[43][1] , \i_fifo_rx/mem[43][0] ,
         \i_fifo_rx/mem[42][7] , \i_fifo_rx/mem[42][6] ,
         \i_fifo_rx/mem[42][5] , \i_fifo_rx/mem[42][4] ,
         \i_fifo_rx/mem[42][3] , \i_fifo_rx/mem[42][2] ,
         \i_fifo_rx/mem[42][1] , \i_fifo_rx/mem[42][0] ,
         \i_fifo_rx/mem[41][7] , \i_fifo_rx/mem[41][6] ,
         \i_fifo_rx/mem[41][5] , \i_fifo_rx/mem[41][4] ,
         \i_fifo_rx/mem[41][3] , \i_fifo_rx/mem[41][2] ,
         \i_fifo_rx/mem[41][1] , \i_fifo_rx/mem[41][0] ,
         \i_fifo_rx/mem[40][7] , \i_fifo_rx/mem[40][6] ,
         \i_fifo_rx/mem[40][5] , \i_fifo_rx/mem[40][4] ,
         \i_fifo_rx/mem[40][3] , \i_fifo_rx/mem[40][2] ,
         \i_fifo_rx/mem[40][1] , \i_fifo_rx/mem[40][0] ,
         \i_fifo_rx/mem[39][7] , \i_fifo_rx/mem[39][6] ,
         \i_fifo_rx/mem[39][5] , \i_fifo_rx/mem[39][4] ,
         \i_fifo_rx/mem[39][3] , \i_fifo_rx/mem[39][2] ,
         \i_fifo_rx/mem[39][1] , \i_fifo_rx/mem[39][0] ,
         \i_fifo_rx/mem[38][7] , \i_fifo_rx/mem[38][6] ,
         \i_fifo_rx/mem[38][5] , \i_fifo_rx/mem[38][4] ,
         \i_fifo_rx/mem[38][3] , \i_fifo_rx/mem[38][2] ,
         \i_fifo_rx/mem[38][1] , \i_fifo_rx/mem[38][0] ,
         \i_fifo_rx/mem[37][7] , \i_fifo_rx/mem[37][6] ,
         \i_fifo_rx/mem[37][5] , \i_fifo_rx/mem[37][4] ,
         \i_fifo_rx/mem[37][3] , \i_fifo_rx/mem[37][2] ,
         \i_fifo_rx/mem[37][1] , \i_fifo_rx/mem[37][0] ,
         \i_fifo_rx/mem[36][7] , \i_fifo_rx/mem[36][6] ,
         \i_fifo_rx/mem[36][5] , \i_fifo_rx/mem[36][4] ,
         \i_fifo_rx/mem[36][3] , \i_fifo_rx/mem[36][2] ,
         \i_fifo_rx/mem[36][1] , \i_fifo_rx/mem[36][0] ,
         \i_fifo_rx/mem[35][7] , \i_fifo_rx/mem[35][6] ,
         \i_fifo_rx/mem[35][5] , \i_fifo_rx/mem[35][4] ,
         \i_fifo_rx/mem[35][3] , \i_fifo_rx/mem[35][2] ,
         \i_fifo_rx/mem[35][1] , \i_fifo_rx/mem[35][0] ,
         \i_fifo_rx/mem[34][7] , \i_fifo_rx/mem[34][6] ,
         \i_fifo_rx/mem[34][5] , \i_fifo_rx/mem[34][4] ,
         \i_fifo_rx/mem[34][3] , \i_fifo_rx/mem[34][2] ,
         \i_fifo_rx/mem[34][1] , \i_fifo_rx/mem[34][0] ,
         \i_fifo_rx/mem[33][7] , \i_fifo_rx/mem[33][6] ,
         \i_fifo_rx/mem[33][5] , \i_fifo_rx/mem[33][4] ,
         \i_fifo_rx/mem[33][3] , \i_fifo_rx/mem[33][2] ,
         \i_fifo_rx/mem[33][1] , \i_fifo_rx/mem[33][0] ,
         \i_fifo_rx/mem[32][7] , \i_fifo_rx/mem[32][6] ,
         \i_fifo_rx/mem[32][5] , \i_fifo_rx/mem[32][4] ,
         \i_fifo_rx/mem[32][3] , \i_fifo_rx/mem[32][2] ,
         \i_fifo_rx/mem[32][1] , \i_fifo_rx/mem[32][0] ,
         \i_fifo_rx/mem[31][7] , \i_fifo_rx/mem[31][6] ,
         \i_fifo_rx/mem[31][5] , \i_fifo_rx/mem[31][4] ,
         \i_fifo_rx/mem[31][3] , \i_fifo_rx/mem[31][2] ,
         \i_fifo_rx/mem[31][1] , \i_fifo_rx/mem[31][0] ,
         \i_fifo_rx/mem[30][7] , \i_fifo_rx/mem[30][6] ,
         \i_fifo_rx/mem[30][5] , \i_fifo_rx/mem[30][4] ,
         \i_fifo_rx/mem[30][3] , \i_fifo_rx/mem[30][2] ,
         \i_fifo_rx/mem[30][1] , \i_fifo_rx/mem[30][0] ,
         \i_fifo_rx/mem[29][7] , \i_fifo_rx/mem[29][6] ,
         \i_fifo_rx/mem[29][5] , \i_fifo_rx/mem[29][4] ,
         \i_fifo_rx/mem[29][3] , \i_fifo_rx/mem[29][2] ,
         \i_fifo_rx/mem[29][1] , \i_fifo_rx/mem[29][0] ,
         \i_fifo_rx/mem[28][7] , \i_fifo_rx/mem[28][6] ,
         \i_fifo_rx/mem[28][5] , \i_fifo_rx/mem[28][4] ,
         \i_fifo_rx/mem[28][3] , \i_fifo_rx/mem[28][2] ,
         \i_fifo_rx/mem[28][1] , \i_fifo_rx/mem[28][0] ,
         \i_fifo_rx/mem[27][7] , \i_fifo_rx/mem[27][6] ,
         \i_fifo_rx/mem[27][5] , \i_fifo_rx/mem[27][4] ,
         \i_fifo_rx/mem[27][3] , \i_fifo_rx/mem[27][2] ,
         \i_fifo_rx/mem[27][1] , \i_fifo_rx/mem[27][0] ,
         \i_fifo_rx/mem[26][7] , \i_fifo_rx/mem[26][6] ,
         \i_fifo_rx/mem[26][5] , \i_fifo_rx/mem[26][4] ,
         \i_fifo_rx/mem[26][3] , \i_fifo_rx/mem[26][2] ,
         \i_fifo_rx/mem[26][1] , \i_fifo_rx/mem[26][0] ,
         \i_fifo_rx/mem[25][7] , \i_fifo_rx/mem[25][6] ,
         \i_fifo_rx/mem[25][5] , \i_fifo_rx/mem[25][4] ,
         \i_fifo_rx/mem[25][3] , \i_fifo_rx/mem[25][2] ,
         \i_fifo_rx/mem[25][1] , \i_fifo_rx/mem[25][0] ,
         \i_fifo_rx/mem[24][7] , \i_fifo_rx/mem[24][6] ,
         \i_fifo_rx/mem[24][5] , \i_fifo_rx/mem[24][4] ,
         \i_fifo_rx/mem[24][3] , \i_fifo_rx/mem[24][2] ,
         \i_fifo_rx/mem[24][1] , \i_fifo_rx/mem[24][0] ,
         \i_fifo_rx/mem[23][7] , \i_fifo_rx/mem[23][6] ,
         \i_fifo_rx/mem[23][5] , \i_fifo_rx/mem[23][4] ,
         \i_fifo_rx/mem[23][3] , \i_fifo_rx/mem[23][2] ,
         \i_fifo_rx/mem[23][1] , \i_fifo_rx/mem[23][0] ,
         \i_fifo_rx/mem[22][7] , \i_fifo_rx/mem[22][6] ,
         \i_fifo_rx/mem[22][5] , \i_fifo_rx/mem[22][4] ,
         \i_fifo_rx/mem[22][3] , \i_fifo_rx/mem[22][2] ,
         \i_fifo_rx/mem[22][1] , \i_fifo_rx/mem[22][0] ,
         \i_fifo_rx/mem[21][7] , \i_fifo_rx/mem[21][6] ,
         \i_fifo_rx/mem[21][5] , \i_fifo_rx/mem[21][4] ,
         \i_fifo_rx/mem[21][3] , \i_fifo_rx/mem[21][2] ,
         \i_fifo_rx/mem[21][1] , \i_fifo_rx/mem[21][0] ,
         \i_fifo_rx/mem[20][7] , \i_fifo_rx/mem[20][6] ,
         \i_fifo_rx/mem[20][5] , \i_fifo_rx/mem[20][4] ,
         \i_fifo_rx/mem[20][3] , \i_fifo_rx/mem[20][2] ,
         \i_fifo_rx/mem[20][1] , \i_fifo_rx/mem[20][0] ,
         \i_fifo_rx/mem[19][7] , \i_fifo_rx/mem[19][6] ,
         \i_fifo_rx/mem[19][5] , \i_fifo_rx/mem[19][4] ,
         \i_fifo_rx/mem[19][3] , \i_fifo_rx/mem[19][2] ,
         \i_fifo_rx/mem[19][1] , \i_fifo_rx/mem[19][0] ,
         \i_fifo_rx/mem[18][7] , \i_fifo_rx/mem[18][6] ,
         \i_fifo_rx/mem[18][5] , \i_fifo_rx/mem[18][4] ,
         \i_fifo_rx/mem[18][3] , \i_fifo_rx/mem[18][2] ,
         \i_fifo_rx/mem[18][1] , \i_fifo_rx/mem[18][0] ,
         \i_fifo_rx/mem[17][7] , \i_fifo_rx/mem[17][6] ,
         \i_fifo_rx/mem[17][5] , \i_fifo_rx/mem[17][4] ,
         \i_fifo_rx/mem[17][3] , \i_fifo_rx/mem[17][2] ,
         \i_fifo_rx/mem[17][1] , \i_fifo_rx/mem[17][0] ,
         \i_fifo_rx/mem[16][7] , \i_fifo_rx/mem[16][6] ,
         \i_fifo_rx/mem[16][5] , \i_fifo_rx/mem[16][4] ,
         \i_fifo_rx/mem[16][3] , \i_fifo_rx/mem[16][2] ,
         \i_fifo_rx/mem[16][1] , \i_fifo_rx/mem[16][0] ,
         \i_fifo_rx/mem[15][7] , \i_fifo_rx/mem[15][6] ,
         \i_fifo_rx/mem[15][5] , \i_fifo_rx/mem[15][4] ,
         \i_fifo_rx/mem[15][3] , \i_fifo_rx/mem[15][2] ,
         \i_fifo_rx/mem[15][1] , \i_fifo_rx/mem[15][0] ,
         \i_fifo_rx/mem[14][7] , \i_fifo_rx/mem[14][6] ,
         \i_fifo_rx/mem[14][5] , \i_fifo_rx/mem[14][4] ,
         \i_fifo_rx/mem[14][3] , \i_fifo_rx/mem[14][2] ,
         \i_fifo_rx/mem[14][1] , \i_fifo_rx/mem[14][0] ,
         \i_fifo_rx/mem[13][7] , \i_fifo_rx/mem[13][6] ,
         \i_fifo_rx/mem[13][5] , \i_fifo_rx/mem[13][4] ,
         \i_fifo_rx/mem[13][3] , \i_fifo_rx/mem[13][2] ,
         \i_fifo_rx/mem[13][1] , \i_fifo_rx/mem[13][0] ,
         \i_fifo_rx/mem[12][7] , \i_fifo_rx/mem[12][6] ,
         \i_fifo_rx/mem[12][5] , \i_fifo_rx/mem[12][4] ,
         \i_fifo_rx/mem[12][3] , \i_fifo_rx/mem[12][2] ,
         \i_fifo_rx/mem[12][1] , \i_fifo_rx/mem[12][0] ,
         \i_fifo_rx/mem[11][7] , \i_fifo_rx/mem[11][6] ,
         \i_fifo_rx/mem[11][5] , \i_fifo_rx/mem[11][4] ,
         \i_fifo_rx/mem[11][3] , \i_fifo_rx/mem[11][2] ,
         \i_fifo_rx/mem[11][1] , \i_fifo_rx/mem[11][0] ,
         \i_fifo_rx/mem[10][7] , \i_fifo_rx/mem[10][6] ,
         \i_fifo_rx/mem[10][5] , \i_fifo_rx/mem[10][4] ,
         \i_fifo_rx/mem[10][3] , \i_fifo_rx/mem[10][2] ,
         \i_fifo_rx/mem[10][1] , \i_fifo_rx/mem[10][0] , \i_fifo_rx/mem[9][7] ,
         \i_fifo_rx/mem[9][6] , \i_fifo_rx/mem[9][5] , \i_fifo_rx/mem[9][4] ,
         \i_fifo_rx/mem[9][3] , \i_fifo_rx/mem[9][2] , \i_fifo_rx/mem[9][1] ,
         \i_fifo_rx/mem[9][0] , \i_fifo_rx/mem[8][7] , \i_fifo_rx/mem[8][6] ,
         \i_fifo_rx/mem[8][5] , \i_fifo_rx/mem[8][4] , \i_fifo_rx/mem[8][3] ,
         \i_fifo_rx/mem[8][2] , \i_fifo_rx/mem[8][1] , \i_fifo_rx/mem[8][0] ,
         \i_fifo_rx/mem[7][7] , \i_fifo_rx/mem[7][6] , \i_fifo_rx/mem[7][5] ,
         \i_fifo_rx/mem[7][4] , \i_fifo_rx/mem[7][3] , \i_fifo_rx/mem[7][2] ,
         \i_fifo_rx/mem[7][1] , \i_fifo_rx/mem[7][0] , \i_fifo_rx/mem[6][7] ,
         \i_fifo_rx/mem[6][6] , \i_fifo_rx/mem[6][5] , \i_fifo_rx/mem[6][4] ,
         \i_fifo_rx/mem[6][3] , \i_fifo_rx/mem[6][2] , \i_fifo_rx/mem[6][1] ,
         \i_fifo_rx/mem[6][0] , \i_fifo_rx/mem[5][7] , \i_fifo_rx/mem[5][6] ,
         \i_fifo_rx/mem[5][5] , \i_fifo_rx/mem[5][4] , \i_fifo_rx/mem[5][3] ,
         \i_fifo_rx/mem[5][2] , \i_fifo_rx/mem[5][1] , \i_fifo_rx/mem[5][0] ,
         \i_fifo_rx/mem[4][7] , \i_fifo_rx/mem[4][6] , \i_fifo_rx/mem[4][5] ,
         \i_fifo_rx/mem[4][4] , \i_fifo_rx/mem[4][3] , \i_fifo_rx/mem[4][2] ,
         \i_fifo_rx/mem[4][1] , \i_fifo_rx/mem[4][0] , \i_fifo_rx/mem[3][7] ,
         \i_fifo_rx/mem[3][6] , \i_fifo_rx/mem[3][5] , \i_fifo_rx/mem[3][4] ,
         \i_fifo_rx/mem[3][3] , \i_fifo_rx/mem[3][2] , \i_fifo_rx/mem[3][1] ,
         \i_fifo_rx/mem[3][0] , \i_fifo_rx/mem[2][7] , \i_fifo_rx/mem[2][6] ,
         \i_fifo_rx/mem[2][5] , \i_fifo_rx/mem[2][4] , \i_fifo_rx/mem[2][3] ,
         \i_fifo_rx/mem[2][2] , \i_fifo_rx/mem[2][1] , \i_fifo_rx/mem[2][0] ,
         \i_fifo_rx/mem[1][7] , \i_fifo_rx/mem[1][6] , \i_fifo_rx/mem[1][5] ,
         \i_fifo_rx/mem[1][4] , \i_fifo_rx/mem[1][3] , \i_fifo_rx/mem[1][2] ,
         \i_fifo_rx/mem[1][1] , \i_fifo_rx/mem[1][0] , \i_fifo_rx/mem[0][7] ,
         \i_fifo_rx/mem[0][6] , \i_fifo_rx/mem[0][5] , \i_fifo_rx/mem[0][4] ,
         \i_fifo_rx/mem[0][3] , \i_fifo_rx/mem[0][2] , \i_fifo_rx/mem[0][1] ,
         \i_fifo_rx/mem[0][0] , \i_fifo_rx/N68 , \i_fifo_rx/N67 ,
         \i_fifo_rx/N66 , \i_fifo_rx/N65 , \i_fifo_rx/N64 , \i_fifo_rx/N63 ,
         \i_fifo_rx/N62 , \i_fifo_rx/N61 , \i_fifo_rx/N59 , \i_fifo_rx/N58 ,
         \i_fifo_rx/N57 , \i_fifo_rx/N56 , \i_fifo_rx/N55 , \i_fifo_rx/N54 ,
         \i_fifo_rx/N46 , \i_fifo_rx/rd_ptr[6] , \i_fifo_rx/wr_ptr[6] ,
         \i_fifo_rx/N44 , \i_fifo_rx/N43 , \i_fifo_rx/N42 , \i_fifo_rx/N41 ,
         \i_fifo_rx/N40 , \i_fifo_rx/N39 , \i_fifo_rx/N38 , \i_fifo_rx/N37 ,
         \i_fifo_rx/N36 , \i_fifo_rx/N35 , \i_mod_iq/fsm_mapping/n232 ,
         \i_mod_iq/fsm_mapping/n231 , \i_mod_iq/fsm_mapping/n230 ,
         \i_mod_iq/fsm_mapping/n229 , \i_mod_iq/fsm_mapping/n228 ,
         \i_mod_iq/fsm_mapping/n227 , \i_mod_iq/fsm_mapping/n226 ,
         \i_mod_iq/fsm_mapping/n225 , \i_mod_iq/fsm_mapping/n224 ,
         \i_mod_iq/fsm_mapping/n223 , \i_mod_iq/fsm_mapping/n222 ,
         \i_mod_iq/fsm_mapping/n221 , \i_mod_iq/fsm_mapping/n220 ,
         \i_mod_iq/fsm_mapping/n218 , \i_mod_iq/fsm_mapping/n217 ,
         \i_mod_iq/fsm_mapping/n216 , \i_mod_iq/fsm_mapping/n215 ,
         \i_mod_iq/fsm_mapping/n214 , \i_mod_iq/fsm_mapping/n213 ,
         \i_mod_iq/fsm_mapping/n212 , \i_mod_iq/fsm_mapping/n211 ,
         \i_mod_iq/fsm_mapping/n210 , \i_mod_iq/fsm_mapping/n209 ,
         \i_mod_iq/fsm_mapping/n208 , \i_mod_iq/fsm_mapping/n207 ,
         \i_mod_iq/fsm_mapping/n206 , \i_mod_iq/fsm_mapping/n205 ,
         \i_mod_iq/fsm_mapping/n204 , \i_mod_iq/fsm_mapping/n203 ,
         \i_mod_iq/fsm_mapping/n202 , \i_mod_iq/fsm_mapping/n201 ,
         \i_mod_iq/fsm_mapping/n199 , \i_mod_iq/fsm_mapping/n197 ,
         \i_mod_iq/fsm_mapping/n196 , \i_mod_iq/fsm_mapping/n195 ,
         \i_mod_iq/fsm_mapping/n194 , \i_mod_iq/fsm_mapping/n193 ,
         \i_mod_iq/fsm_mapping/n192 , \i_mod_iq/fsm_mapping/n191 ,
         \i_mod_iq/fsm_mapping/n188 , \i_mod_iq/fsm_mapping/n187 ,
         \i_mod_iq/fsm_mapping/n185 , \i_mod_iq/fsm_mapping/n184 ,
         \i_mod_iq/fsm_mapping/n183 , \i_mod_iq/fsm_mapping/n182 ,
         \i_mod_iq/fsm_mapping/n181 , \i_mod_iq/fsm_mapping/n180 ,
         \i_mod_iq/fsm_mapping/n179 , \i_mod_iq/fsm_mapping/n178 ,
         \i_mod_iq/fsm_mapping/n177 , \i_mod_iq/fsm_mapping/n175 ,
         \i_mod_iq/fsm_mapping/n174 , \i_mod_iq/fsm_mapping/n173 ,
         \i_mod_iq/fsm_mapping/n171 , \i_mod_iq/fsm_mapping/n170 ,
         \i_mod_iq/fsm_mapping/n169 , \i_mod_iq/fsm_mapping/n168 ,
         \i_mod_iq/fsm_mapping/n167 , \i_mod_iq/fsm_mapping/n166 ,
         \i_mod_iq/fsm_mapping/n165 , \i_mod_iq/fsm_mapping/n164 ,
         \i_mod_iq/fsm_mapping/n163 , \i_mod_iq/fsm_mapping/n161 ,
         \i_mod_iq/fsm_mapping/n160 , \i_mod_iq/fsm_mapping/n159 ,
         \i_mod_iq/fsm_mapping/n158 , \i_mod_iq/fsm_mapping/n157 ,
         \i_mod_iq/fsm_mapping/n156 , \i_mod_iq/fsm_mapping/n155 ,
         \i_mod_iq/fsm_mapping/n154 , \i_mod_iq/fsm_mapping/n153 ,
         \i_mod_iq/fsm_mapping/n152 , \i_mod_iq/fsm_mapping/n151 ,
         \i_mod_iq/fsm_mapping/n150 , \i_mod_iq/fsm_mapping/n149 ,
         \i_mod_iq/fsm_mapping/n148 , \i_mod_iq/fsm_mapping/n147 ,
         \i_mod_iq/fsm_mapping/n146 , \i_mod_iq/fsm_mapping/n145 ,
         \i_mod_iq/fsm_mapping/n143 , \i_mod_iq/fsm_mapping/n140 ,
         \i_mod_iq/fsm_mapping/n139 , \i_mod_iq/fsm_mapping/n138 ,
         \i_mod_iq/fsm_mapping/n137 , \i_mod_iq/fsm_mapping/n136 ,
         \i_mod_iq/fsm_mapping/n135 , \i_mod_iq/fsm_mapping/n134 ,
         \i_mod_iq/fsm_mapping/n133 , \i_mod_iq/fsm_mapping/n132 ,
         \i_mod_iq/fsm_mapping/n131 , \i_mod_iq/fsm_mapping/n130 ,
         \i_mod_iq/fsm_mapping/n129 , \i_mod_iq/fsm_mapping/n128 ,
         \i_mod_iq/fsm_mapping/n127 , \i_mod_iq/fsm_mapping/n126 ,
         \i_mod_iq/fsm_mapping/n125 , \i_mod_iq/fsm_mapping/n124 ,
         \i_mod_iq/fsm_mapping/n123 , \i_mod_iq/fsm_mapping/n120 ,
         \i_mod_iq/fsm_mapping/n119 , \i_mod_iq/fsm_mapping/n118 ,
         \i_mod_iq/fsm_mapping/n117 , \i_mod_iq/fsm_mapping/n116 ,
         \i_mod_iq/fsm_mapping/n115 , \i_mod_iq/fsm_mapping/n114 ,
         \i_mod_iq/fsm_mapping/n113 , \i_mod_iq/fsm_mapping/n112 ,
         \i_mod_iq/fsm_mapping/n111 , \i_mod_iq/fsm_mapping/n110 ,
         \i_mod_iq/fsm_mapping/n109 , \i_mod_iq/fsm_mapping/n108 ,
         \i_mod_iq/fsm_mapping/n107 , \i_mod_iq/fsm_mapping/n106 ,
         \i_mod_iq/fsm_mapping/n105 , \i_mod_iq/fsm_mapping/n104 ,
         \i_mod_iq/fsm_mapping/n103 , \i_mod_iq/fsm_mapping/n102 ,
         \i_mod_iq/fsm_mapping/n101 , \i_mod_iq/fsm_mapping/n100 ,
         \i_mod_iq/fsm_mapping/n99 , \i_mod_iq/fsm_mapping/n98 ,
         \i_mod_iq/fsm_mapping/n97 , \i_mod_iq/fsm_mapping/n96 ,
         \i_mod_iq/fsm_mapping/n95 , \i_mod_iq/fsm_mapping/n94 ,
         \i_mod_iq/fsm_mapping/n93 , \i_mod_iq/fsm_mapping/n92 ,
         \i_mod_iq/fsm_mapping/n90 , \i_mod_iq/fsm_mapping/n89 ,
         \i_mod_iq/fsm_mapping/n88 , \i_mod_iq/fsm_mapping/n87 ,
         \i_mod_iq/fsm_mapping/n86 , \i_mod_iq/fsm_mapping/n85 ,
         \i_mod_iq/fsm_mapping/n84 , \i_mod_iq/fsm_mapping/n83 ,
         \i_mod_iq/fsm_mapping/n82 , \i_mod_iq/fsm_mapping/n81 ,
         \i_mod_iq/fsm_mapping/n80 , \i_mod_iq/fsm_mapping/n79 ,
         \i_mod_iq/fsm_mapping/n77 , \i_mod_iq/fsm_mapping/n76 ,
         \i_mod_iq/fsm_mapping/n75 , \i_mod_iq/fsm_mapping/n74 ,
         \i_mod_iq/fsm_mapping/n73 , \i_mod_iq/fsm_mapping/n72 ,
         \i_mod_iq/fsm_mapping/n71 , \i_mod_iq/fsm_mapping/n70 ,
         \i_mod_iq/fsm_mapping/n69 , \i_mod_iq/fsm_mapping/n68 ,
         \i_mod_iq/fsm_mapping/n67 , \i_mod_iq/fsm_mapping/n66 ,
         \i_mod_iq/fsm_mapping/n65 , \i_mod_iq/fsm_mapping/n64 ,
         \i_mod_iq/fsm_mapping/n63 , \i_mod_iq/fsm_mapping/n62 ,
         \i_mod_iq/fsm_mapping/n61 , \i_mod_iq/fsm_mapping/n60 ,
         \i_mod_iq/fsm_mapping/n59 , \i_mod_iq/fsm_mapping/n58 ,
         \i_mod_iq/fsm_mapping/n57 , \i_mod_iq/fsm_mapping/n56 ,
         \i_mod_iq/fsm_mapping/n55 , \i_mod_iq/fsm_mapping/n54 ,
         \i_mod_iq/fsm_mapping/n53 , \i_mod_iq/fsm_mapping/n52 ,
         \i_mod_iq/fsm_mapping/n51 , \i_mod_iq/fsm_mapping/n50 ,
         \i_mod_iq/fsm_mapping/n49 , \i_mod_iq/fsm_mapping/n48 ,
         \i_mod_iq/fsm_mapping/n47 , \i_mod_iq/fsm_mapping/n46 ,
         \i_mod_iq/fsm_mapping/n45 , \i_mod_iq/fsm_mapping/n44 ,
         \i_mod_iq/fsm_mapping/n43 , \i_mod_iq/fsm_mapping/n42 ,
         \i_mod_iq/fsm_mapping/n41 , \i_mod_iq/fsm_mapping/n40 ,
         \i_mod_iq/fsm_mapping/n39 , \i_mod_iq/fsm_mapping/n38 ,
         \i_mod_iq/fsm_mapping/n37 , \i_mod_iq/fsm_mapping/n36 ,
         \i_mod_iq/fsm_mapping/n35 , \i_mod_iq/fsm_mapping/n34 ,
         \i_mod_iq/fsm_mapping/n33 , \i_mod_iq/fsm_mapping/n32 ,
         \i_mod_iq/fsm_mapping/n31 , \i_mod_iq/fsm_mapping/n30 ,
         \i_mod_iq/fsm_mapping/n29 , \i_mod_iq/fsm_mapping/n28 ,
         \i_mod_iq/fsm_mapping/N261 , \i_mod_iq/fsm_mapping/N260 ,
         \i_mod_iq/fsm_mapping/N259 , \i_mod_iq/fsm_mapping/s_b_in_prev ,
         \i_mod_iq/fsm_mapping/b_in_prev , \i_mod_iq/fsm_mapping/S_AQ ,
         \i_mod_iq/fsm_mapping/S_AI , \i_mod_iq/fsm_mapping/en_prev ,
         \i_mod_iq/fsm_mapping/en_10MHz_prev , \i_mod_iq/en_gen_map/n4 ,
         \i_mod_iq/en_gen_map/n3 , \i_mod_iq/en_gen_map/n1 ,
         \i_mod_iq/en_gen_map/N13 , \i_mod_iq/en_gen_map/N6 ,
         \i_iq_demod/demod/n43 , \i_iq_demod/demod/n41 ,
         \i_iq_demod/demod/n39 , \i_iq_demod/demod/n37 ,
         \i_iq_demod/demod/n35 , \i_iq_demod/demod/n33 ,
         \i_iq_demod/demod/n32 , \i_iq_demod/demod/n31 ,
         \i_iq_demod/demod/n29 , \i_iq_demod/demod/n27 ,
         \i_iq_demod/demod/n25 , \i_iq_demod/demod/n23 ,
         \i_iq_demod/demod/n22 , \i_iq_demod/demod/n20 ,
         \i_iq_demod/demod/dp_cluster_1/N85 ,
         \i_iq_demod/demod/dp_cluster_1/N86 ,
         \i_iq_demod/demod/dp_cluster_1/N87 ,
         \i_iq_demod/demod/dp_cluster_1/N88 ,
         \i_iq_demod/demod/dp_cluster_0/N90 ,
         \i_iq_demod/demod/dp_cluster_0/N91 ,
         \i_iq_demod/demod/dp_cluster_0/N92 ,
         \i_iq_demod/demod/dp_cluster_0/N93 , \i_iq_demod/demod/N41 ,
         \i_iq_demod/demod/N36 , \i_iq_demod/filtre_I/n42 ,
         \i_iq_demod/filtre_I/n22 , \i_iq_demod/filtre_I/n10 ,
         \i_iq_demod/filtre_I/n9 , \i_iq_demod/filtre_I/n7 ,
         \i_iq_demod/filtre_I/n6 , \i_iq_demod/filtre_I/n4 ,
         \i_iq_demod/filtre_I/n2 , \i_iq_demod/filtre_I/n1 ,
         \i_iq_demod/filtre_I/N123 , \i_iq_demod/filtre_I/_16_net_[8] ,
         \i_iq_demod/filtre_I/_15_net_[8] , \i_iq_demod/filtre_I/N28 ,
         \i_iq_demod/filtre_I/N27 , \i_iq_demod/filtre_I/N26 ,
         \i_iq_demod/filtre_I/N25 , \i_iq_demod/filtre_I/N24 ,
         \i_iq_demod/filtre_I/N23 , \i_iq_demod/filtre_I/N22 ,
         \i_iq_demod/filtre_I/N21 , \i_iq_demod/filtre_I/N20 ,
         \i_iq_demod/filtre_I/N19 , \i_iq_demod/filtre_I/N18 ,
         \i_iq_demod/filtre_I/N17 , \i_iq_demod/filtre_I/N16 ,
         \i_iq_demod/filtre_I/N15 , \i_iq_demod/gen_sin/n22 ,
         \i_iq_demod/gen_sin/n21 , \i_iq_demod/gen_sin/n20 ,
         \i_iq_demod/gen_sin/n19 , \i_iq_demod/gen_sin/n18 ,
         \i_iq_demod/gen_sin/n6 , \i_iq_demod/gen_sin/n5 ,
         \i_iq_demod/gen_sin/n3 , \i_iq_demod/gen_sin/n2 ,
         \i_iq_demod/gen_sin/n1 , \i_iq_demod/gen_sin/N106 ,
         \i_iq_demod/gen_sin/N17 , \i_iq_demod/gen_sin/N15 , \i_cordic/S0/n39 ,
         \i_cordic/S0/n37 , \i_cordic/S0/n35 , \i_cordic/S0/n34 ,
         \i_cordic/S0/n33 , \i_cordic/S0/n29 , \i_cordic/S0/n28 ,
         \i_cordic/S0/n27 , \i_cordic/S0/n26 , \i_cordic/S0/n25 ,
         \i_cordic/S0/n24 , \i_cordic/S0/n23 , \i_cordic/S0/n22 ,
         \i_cordic/S0/N32 , \i_cordic/S0/N19 , \i_cordic/S0/N18 ,
         \i_cordic/S0/N17 , \i_cordic/S0/N16 , \i_cordic/S0/N14 ,
         \i_cordic/S0/N13 , \i_cordic/S0/N12 , \i_cordic/S0/N11 ,
         \i_cordic/S0/N10 , \i_cordic/S0/N9 , \i_cordic/S0/N7 ,
         \i_cordic/S0/N6 , \i_cordic/S0/N5 , \i_cordic/S0/N4 ,
         \i_cordic/S1/n35 , \i_cordic/S1/n34 , \i_cordic/S1/N38 ,
         \i_cordic/S1/N26 , \i_cordic/S1/N25 , \i_cordic/S1/N24 ,
         \i_cordic/S1/N23 , \i_cordic/S1/N22 , \i_cordic/S1/N21 ,
         \i_cordic/S1/N20 , \i_cordic/S1/N19 , \i_cordic/S1/N18 ,
         \i_cordic/S1/N17 , \i_cordic/S1/N16 , \i_cordic/S1/N15 ,
         \i_cordic/S1/N14 , \i_cordic/S1/N13 , \i_cordic/S1/N12 ,
         \i_cordic/S1/N11 , \i_cordic/S1/N8 , \i_cordic/S1/N7 ,
         \i_cordic/S1/N6 , \i_cordic/S1/N5 , \i_cordic/S2/n37 ,
         \i_cordic/S2/n36 , \i_cordic/S2/n35 , \i_cordic/S2/n34 ,
         \i_cordic/S2/n21 , \i_cordic/S2/N38 , \i_cordic/S2/N37 ,
         \i_cordic/S2/N36 , \i_cordic/S2/N32 , \i_cordic/S2/N31 ,
         \i_cordic/S2/N30 , \i_cordic/S2/N29 , \i_cordic/S2/N26 ,
         \i_cordic/S2/N20 , \i_cordic/S3/n30 , \i_cordic/S3/n28 ,
         \i_cordic/S3/N37 , \i_cordic/S3/N36 , \i_cdr/i_bit_recovery/n33 ,
         \i_cdr/i_bit_recovery/n32 , \i_cdr/i_bit_recovery/n31 ,
         \i_cdr/i_bit_recovery/n30 , \i_cdr/i_bit_recovery/n29 ,
         \i_cdr/i_bit_recovery/n28 , \i_cdr/i_bit_recovery/n27 ,
         \i_cdr/i_bit_recovery/n26 , \i_cdr/i_bit_recovery/n25 ,
         \i_cdr/i_bit_recovery/n14 , \i_cdr/i_bit_recovery/n12 ,
         \i_cdr/i_bit_recovery/n11 , \i_cdr/i_bit_recovery/n10 ,
         \i_cdr/i_bit_recovery/n9 , \i_cdr/i_bit_recovery/n8 ,
         \i_cdr/i_bit_recovery/N91 , \i_cdr/i_bit_recovery/phase_diff[5] ,
         \i_cdr/i_cdr/n29 , \i_cdr/i_cdr/n28 , \i_cdr/i_cdr/n27 ,
         \i_cdr/i_cdr/n12 , \i_cdr/i_cdr/n11 , \i_cdr/i_cdr/n9 ,
         \i_cdr/i_cdr/n8 , \i_cdr/i_cdr/n7 , \i_cdr/i_cdr/n6 ,
         \i_cdr/i_cdr/n5 , \i_cdr/i_cdr/n4 , \i_cdr/i_cdr/n3 ,
         \i_cdr/i_cdr/N160 , \i_cdr/i_cdr/N157 , \i_cdr/i_cdr/N156 ,
         \i_cdr/i_cdr/N155 , \i_cdr/i_cdr/N154 , \i_cdr/i_cdr/N153 ,
         \i_cdr/i_cdr/N151 , \i_cdr/i_cdr/N150 , \i_cdr/i_cdr/N149 ,
         \i_cdr/i_cdr/N145 , \i_cdr/i_cdr/cycles[2] ,
         \i_cdr/i_cdr/curr_state[1] , \i_cdr/i_cdr/N17 , \i_cdr/i_cdr/q3 ,
         \i_cdr/i_cdr/data_en_w , \i_cdr/i_cdr/q4 , \i_cdr/i_cdr/q2 ,
         \i_cdr/i_cdr/q1 , \i_iq_demod/demod/validation/n5 ,
         \i_iq_demod/demod/validation/n3 , \i_iq_demod/demod/validation/n2 ,
         \i_iq_demod/demod/validation/n1 , \i_iq_demod/filtre_I/data_reg1/n36 ,
         \i_iq_demod/filtre_I/data_reg1/n35 ,
         \i_iq_demod/filtre_I/data_reg1/n34 ,
         \i_iq_demod/filtre_I/data_reg1/n33 ,
         \i_iq_demod/filtre_I/data_reg1/n32 ,
         \i_iq_demod/filtre_I/data_reg1/n31 ,
         \i_iq_demod/filtre_I/data_reg1/n30 ,
         \i_iq_demod/filtre_I/data_reg1/n29 ,
         \i_iq_demod/filtre_I/data_reg1/n28 ,
         \i_iq_demod/filtre_I/data_reg1/n27 ,
         \i_iq_demod/filtre_I/data_reg1/n26 ,
         \i_iq_demod/filtre_I/data_reg1/n25 ,
         \i_iq_demod/filtre_I/data_reg1/n24 ,
         \i_iq_demod/filtre_I/data_reg1/n23 ,
         \i_iq_demod/filtre_I/data_reg1/n22 ,
         \i_iq_demod/filtre_I/data_reg1/n21 ,
         \i_iq_demod/filtre_I/data_reg1/n20 ,
         \i_iq_demod/filtre_I/data_reg1/n19 ,
         \i_iq_demod/filtre_I/data_reg1/n18 ,
         \i_iq_demod/filtre_I/data_reg1/n17 ,
         \i_iq_demod/filtre_I/data_reg1/n16 ,
         \i_iq_demod/filtre_I/data_reg1/n15 ,
         \i_iq_demod/filtre_I/data_reg1/n14 ,
         \i_iq_demod/filtre_I/data_reg1/n13 ,
         \i_iq_demod/filtre_I/data_reg1/n12 ,
         \i_iq_demod/filtre_I/data_reg1/n11 ,
         \i_iq_demod/filtre_I/data_reg1/n10 ,
         \i_iq_demod/filtre_I/data_reg1/n9 ,
         \i_iq_demod/filtre_I/data_reg1/n8 ,
         \i_iq_demod/filtre_I/data_reg1/n7 ,
         \i_iq_demod/filtre_I/data_reg1/n6 ,
         \i_iq_demod/filtre_I/data_reg1/n5 ,
         \i_iq_demod/filtre_I/data_reg1/n4 ,
         \i_iq_demod/filtre_I/data_reg1/n3 ,
         \i_iq_demod/filtre_I/data_reg1/n2 ,
         \i_iq_demod/filtre_I/data_reg1/n1 , \i_iq_demod/filtre_I/factor/n57 ,
         \i_iq_demod/filtre_I/factor/n52 , \i_iq_demod/filtre_I/factor/n42 ,
         \i_iq_demod/filtre_I/factor/n39 , \i_iq_demod/filtre_I/factor/n26 ,
         \i_iq_demod/filtre_I/factor/n24 , \i_iq_demod/filtre_I/factor/n23 ,
         \i_iq_demod/filtre_I/factor/n11 , \i_iq_demod/filtre_I/factor/n8 ,
         \i_iq_demod/filtre_I/factor/n7 , \i_iq_demod/filtre_I/factor/n6 ,
         \i_iq_demod/filtre_I/factor/n5 , \i_iq_demod/filtre_I/factor/n4 ,
         \i_iq_demod/filtre_I/shift_r/n6 , \i_iq_demod/filtre_I/shift_r/n5 ,
         \i_iq_demod/filtre_I/shift_r/n3 , \i_iq_demod/filtre_I/shift_r/n2 ,
         \i_iq_demod/filtre_I/shift_r/n1 , \i_iq_demod/filtre_I/shift_r/N9 ,
         \i_iq_demod/filtre_I/shift_r/N8 , \i_iq_demod/filtre_I/shift_r/N3 ,
         \i_iq_demod/filtre_I/temp_adder/n57 ,
         \i_iq_demod/filtre_I/temp_adder/n54 ,
         \i_iq_demod/filtre_I/temp_adder/n51 ,
         \i_iq_demod/filtre_I/temp_adder/n48 ,
         \i_iq_demod/filtre_I/temp_adder/n45 ,
         \i_iq_demod/filtre_I/temp_adder/n42 ,
         \i_iq_demod/filtre_I/temp_adder/n41 ,
         \i_iq_demod/filtre_I/temp_adder/n40 ,
         \i_iq_demod/filtre_I/temp_adder/n38 ,
         \i_iq_demod/filtre_I/temp_adder/n35 ,
         \i_iq_demod/filtre_I/temp_adder/n33 ,
         \i_iq_demod/filtre_I/temp_adder/n20 ,
         \i_iq_demod/filtre_I/temp_adder/n18 ,
         \i_iq_demod/filtre_I/temp_adder/n17 ,
         \i_iq_demod/filtre_I/temp_adder/n15 ,
         \i_iq_demod/filtre_I/temp_adder/n14 ,
         \i_iq_demod/filtre_I/temp_adder/n13 ,
         \i_iq_demod/filtre_I/temp_adder/n11 ,
         \i_iq_demod/filtre_I/temp_adder/n10 ,
         \i_iq_demod/filtre_I/temp_adder/n9 ,
         \i_iq_demod/filtre_I/temp_adder/n7 ,
         \i_iq_demod/filtre_I/temp_adder/n6 ,
         \i_iq_demod/filtre_I/temp_adder/n5 ,
         \i_iq_demod/filtre_I/temp_adder/n3 ,
         \i_iq_demod/filtre_I/temp_adder/n2 ,
         \i_iq_demod/filtre_I/temp_adder/n1 ,
         \i_iq_demod/filtre_I/sum1_adder/n15 ,
         \i_iq_demod/filtre_I/sum1_adder/n14 ,
         \i_iq_demod/filtre_I/sum1_adder/n7 ,
         \i_iq_demod/filtre_I/sum1_adder/n6 ,
         \i_iq_demod/filtre_I/sum1_adder/n5 ,
         \i_iq_demod/filtre_I/sum1_adder/n4 ,
         \i_iq_demod/filtre_I/mult1_multiplier/n25 ,
         \i_iq_demod/filtre_I/mult1_multiplier/n21 ,
         \i_iq_demod/filtre_I/mult1_multiplier/n20 ,
         \i_iq_demod/filtre_I/mult1_multiplier/n19 ,
         \i_iq_demod/filtre_I/mult1_multiplier/n18 ,
         \i_iq_demod/filtre_I/mult1_multiplier/n17 ,
         \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[9] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[5] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[9] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[5] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[9] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[5] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[9] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[5] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[9] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[5] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/B_pipe ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[12][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[11][1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[11][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[1][6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[1][7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[2][1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[2][3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[2][5] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[2][7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[2][8] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[3][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[3][1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[3][4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[3][5] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[3][6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[3][7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[3][8] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[4][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[4][1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[4][2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[4][3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[4][4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[4][7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[4][8] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[5][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[5][1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[5][2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[5][6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[5][7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[5][8] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[6][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[6][1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[6][2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[6][3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[6][4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[6][7] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[7][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[7][1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[7][2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[7][3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[7][6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[8][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[8][1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[8][2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[8][3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[8][4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[9][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[9][1] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[9][2] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[9][3] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[9][4] ,
         \i_iq_demod/filtre_I/tot_adder/n50 ,
         \i_iq_demod/filtre_I/tot_adder/n39 ,
         \i_iq_demod/filtre_I/tot_adder/n38 ,
         \i_iq_demod/filtre_I/tot_adder/n35 ,
         \i_iq_demod/filtre_I/tot_adder/n34 ,
         \i_iq_demod/filtre_I/tot_adder/n33 ,
         \i_iq_demod/filtre_I/tot_adder/n32 ,
         \i_iq_demod/filtre_I/tot_adder/n31 ,
         \i_iq_demod/filtre_I/tot_adder/n28 ,
         \i_iq_demod/filtre_I/tot_adder/n27 ,
         \i_iq_demod/filtre_I/tot_adder/n18 ,
         \i_iq_demod/filtre_I/tot_adder/n17 ,
         \i_iq_demod/filtre_I/tot_adder/n15 ,
         \i_iq_demod/filtre_I/tot_adder/n14 ,
         \i_iq_demod/filtre_I/tot_adder/n13 ,
         \i_iq_demod/filtre_I/tot_adder/n11 ,
         \i_iq_demod/filtre_I/tot_adder/n10 ,
         \i_iq_demod/filtre_I/tot_adder/n9 ,
         \i_iq_demod/filtre_I/tot_adder/n7 ,
         \i_iq_demod/filtre_I/tot_adder/n6 ,
         \i_iq_demod/filtre_I/tot_adder/n5 ,
         \i_iq_demod/filtre_I/tot_adder/n3 ,
         \i_iq_demod/filtre_I/tot_adder/n2 ,
         \i_iq_demod/filtre_I/tot_adder/n1 ,
         \i_iq_demod/filtre_I/mult1_multiplier/genblk1[0].adder/n10 ,
         \i_iq_demod/filtre_Q/N123 , \i_iq_demod/filtre_Q/_16_net_[8] ,
         \i_iq_demod/filtre_Q/_15_net_[8] , \i_iq_demod/filtre_Q/N28 ,
         \i_iq_demod/filtre_Q/N27 , \i_iq_demod/filtre_Q/N26 ,
         \i_iq_demod/filtre_Q/N25 , \i_iq_demod/filtre_Q/N24 ,
         \i_iq_demod/filtre_Q/N23 , \i_iq_demod/filtre_Q/N22 ,
         \i_iq_demod/filtre_Q/N21 , \i_iq_demod/filtre_Q/N20 ,
         \i_iq_demod/filtre_Q/N19 , \i_iq_demod/filtre_Q/N18 ,
         \i_iq_demod/filtre_Q/N17 , \i_iq_demod/filtre_Q/N16 ,
         \i_iq_demod/filtre_Q/N15 , \i_iq_demod/filtre_Q/shift_r/N9 ,
         \i_iq_demod/filtre_Q/shift_r/N8 , \i_iq_demod/filtre_Q/shift_r/N3 ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[9] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[9] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[9] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[9] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[9] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/B_pipe ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[12][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[11][1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[11][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[1][6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[1][7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[2][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[2][2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[2][4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[2][5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[2][6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[2][7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[2][8] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[3][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[3][1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[3][2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[3][3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[3][5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[3][6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[3][7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[3][8] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[4][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[4][1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[4][2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[4][3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[4][5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[4][6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[4][7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[4][8] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[5][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[5][1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[5][2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[5][3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[5][4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[5][5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[5][6] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[5][7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[5][8] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[6][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[6][2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[6][3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[6][4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[6][5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[6][7] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[7][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[7][1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[7][2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[7][3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[7][4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[7][5] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[8][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[8][1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[8][2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[8][3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[8][4] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[9][0] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[9][1] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[9][2] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[9][3] ,
         \i_iq_demod/filtre_Q/mult2_multiplier/register[9][4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[9] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[9] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[9] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[9] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[9] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/B_pipe ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[12][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[11][1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[11][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[1][6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[1][7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[2][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[2][1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[2][2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[2][3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[2][4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[2][5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[2][6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[2][7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[2][8] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[3][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[3][1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[3][2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[3][3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[3][4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[3][5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[3][6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[3][7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[3][8] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[4][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[4][1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[4][2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[4][3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[4][4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[4][5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[4][6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[4][7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[4][8] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[5][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[5][1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[5][2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[5][3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[5][4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[5][5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[5][6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[5][7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[5][8] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[6][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[6][1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[6][2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[6][3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[6][5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[6][6] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[6][7] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[7][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[7][1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[7][2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[7][3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[7][5] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[8][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[8][1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[8][2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[8][3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[8][4] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[9][0] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[9][1] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[9][2] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[9][3] ,
         \i_iq_demod/filtre_Q/mult1_multiplier/register[9][4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[7] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[7] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[9] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[7] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[9] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[7] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[9] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[7] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[9] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[7] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[9] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/B_pipe ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[12][0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[11][1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[11][0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[1][6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[1][7] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[2][0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[2][1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[2][2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[2][3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[2][4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[2][5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[2][6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[2][7] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[2][8] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[3][1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[3][2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[3][3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[3][4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[3][5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[3][6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[3][7] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[3][8] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[4][0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[4][1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[4][2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[4][3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[4][4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[4][5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[4][6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[4][7] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[4][8] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[5][0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[5][1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[5][2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[5][3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[5][4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[5][5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[5][6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[5][7] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[6][0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[6][1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[6][2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[6][4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[6][5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[6][6] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[7][0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[7][1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[7][2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[7][4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[7][5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[8][0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[8][1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[8][2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[8][3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[8][4] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[8][5] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[9][0] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[9][1] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[9][2] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[9][3] ,
         \i_iq_demod/filtre_I/mult2_multiplier/register[9][4] ,
         \i_cdr/i_bit_recovery/sub_68/carry[5] , \i_cordic/S2/sub_53/carry[5] ,
         \i_cordic/S2/add_53/carry[5] , \i_cordic/S2/sub_56/carry[5] , n83,
         n84, n85, n86, n87, n88, n89, n90, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n161, n162, n163, n164, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n302, n303, n305, n306, n307, n311,
         n314, n315, n316, n317, n318, n319, n321, n324, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n367, n369, n370, n371, n372, n373, n376, n377, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n396, n398, n400, n402, n403, n404, n405, n407, n408,
         n409, n410, n411, n413, n414, n415, n416, n417, n419, n421, n422,
         n423, n424, n426, n428, n438, n441, n442, n444, n446, n447, n448,
         n449, n450, n451, n455, n457, n458, n459, n460, n461, n462, n463,
         n464, n466, n471, n480, n482, n483, n484, n485, n486, n487, n489,
         n497, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n517, n520, n521, n522, n523, n524, n525, n526, n527,
         n532, n534, n535, n536, n537, n539, n540, n541, n542, n544, n546,
         n547, n548, n549, n550, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n585, n587, n589, n591, n592, n593, n594, n596,
         n597, n598, n599, n600, n602, n603, n605, n606, n608, n610, n612,
         n616, n617, n618, n620, n621, n622, n623, n624, n625, n626, n627,
         n629, n630, n631, n632, n634, n635, n636, n638, n639, n640, n641,
         n643, n644, n645, n646, n647, n648, n650, n651, n652, n653, n654,
         n656, n658, n661, n663, n664, n665, n667, n668, n670, n672, n673,
         n674, n675, n676, n677, n679, n683, n684, n685, n686, n687, n690,
         n691, n692, n693, n695, n696, n697, n698, n699, n700, n701, n704,
         n706, n707, n710, n711, n712, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n725, n726, n727, n729, n730, n731, n732, n734,
         n736, n737, n738, n739, n740, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n775, n777, n779, n781, n782, n783, n784,
         n786, n787, n788, n789, n790, n792, n795, n796, n798, n800, n802,
         n804, n805, n806, n807, n808, n810, n811, n812, n813, n814, n816,
         n818, n819, n820, n821, n823, n824, n825, n826, n827, n828, n830,
         n832, n833, n834, n836, n837, n838, n840, n841, n842, n843, n844,
         n845, n846, n847, n849, n850, n851, n852, n853, n856, n857, n859,
         n860, n861, n862, n863, n864, n865, n866, n868, n870, n873, n874,
         n875, n876, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n890, n896, n899, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n911, n914, n915, n916, n918, n919, n920, n921,
         n923, n925, n926, n927, n928, n929, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n964, n965, n966, n967, n968, n970,
         n971, n972, n973, n975, n977, n978, n979, n981, n982, n985, n987,
         n989, n990, n991, n993, n995, n997, n999, n1001, n1002, n1003, n1004,
         n1006, n1008, n1009, n1010, n1011, n1013, n1015, n1016, n1017, n1020,
         n1025, n1026, n1027, n1029, n1030, n1031, n1032, n1033, n1035, n1037,
         n1041, n1043, n1044, n1047, n1049, n1051, n1052, n1053, n1054, n1055,
         n1056, n1058, n1059, n1060, n1063, n1064, n1066, n1071, n1072, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1082, n1084, n1085, n1086,
         n1088, n1089, n1090, n1091, n1093, n1094, n1095, n1096, n1097, n1098,
         n1100, n1101, n1104, n1105, n1106, n1108, n1110, n1111, n1113, n1115,
         n1117, n1118, n1119, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1156, n1157, n1158,
         n1160, n1161, n1162, n1164, n1165, n1166, n1168, n1169, n1170, n1171,
         n1174, n1175, n1176, n1177, n1178, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1214, n1216, n1217,
         n1218, n1219, n1220, n1221, n1223, n1224, n1225, n1226, n1227, n1228,
         n1230, n1231, n1232, n1234, n1235, n1236, n1238, n1239, n1240, n1242,
         n1243, n1244, n1245, n1246, n1248, n1249, n1250, n1251, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, net41341,
         net41344, net41468, net41482, net41535, net41570, net41781, net41786,
         net41833, net42078, net42210, net42536, net42565, net42758, net42841,
         net42857, net42883, net42978, net43019, net43018, net43044, net43064,
         net43117, net43270, net43436, net43481, n432, n431, n429, n427,
         \i_iq_demod/filtre_I/sum1_adder/n8 ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[2][4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[4] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[3] , net42230, net41996,
         net41398, n496, n493,
         \i_iq_demod/filtre_I/mult1_multiplier/register[5][4] , net42279,
         net42278, net41707, n478, n477, n474, n473, n472, n470, n468,
         \i_iq_demod/filtre_I/mult1_multiplier/register[5][5] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[4][6] ,
         \i_iq_demod/filtre_I/mult1_multiplier/register[4][5] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[3] , net42042,
         net42041, net41794, net41766, n530, n529, n528,
         \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[5] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[5] , n439, n437, n435,
         n433, \i_iq_demod/filtre_I/mult1_multiplier/register[2][0] ,
         \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[2] , n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946;
  wire   [3:0] mod_iq_ibb_o;
  wire   [3:0] mod_iq_qbb_o;
  wire   [4:0] demod_iq_iif_i;
  wire   [4:0] demod_iq_qif_i;
  wire   [4:0] demod_iq_ibb_o;
  wire   [4:0] demod_iq_qbb_o;
  wire   [4:0] cordic_ibb_i;
  wire   [4:0] cordic_qbb_i;
  wire   [5:0] cordic_phase_o;
  wire   [5:0] cdr_phase_i;
  wire   [7:0] fifo_rx_prdata_o;
  wire   [4:0] \i_fifo_tx/counter_clock ;
  wire   [4:0] \i_iq_demod/Q_BB_IN ;
  wire   [4:0] \i_iq_demod/I_BB_IN ;
  wire   [1:0] \i_iq_demod/cosine_IN ;
  wire   [1:0] \i_iq_demod/sine_IN ;
  wire   [4:0] \i_cordic/qbb_ibuff ;
  wire   [4:0] \i_cordic/ibb_ibuff ;
  wire   [7:0] \i_fifo_rx/i ;
  wire   [7:0] \i_fifo_rx/shift_register ;
  wire   [1:0] \i_mod_iq/fsm_mapping/N_STATE ;
  wire   [1:0] \i_mod_iq/fsm_mapping/C_STATE ;
  wire   [3:0] \i_mod_iq/fsm_mapping/temp_QBB ;
  wire   [3:0] \i_mod_iq/fsm_mapping/temp_IBB ;
  wire   [2:0] \i_mod_iq/fsm_mapping/cpt_old ;
  wire   [2:0] \i_mod_iq/fsm_mapping/cpt ;
  wire   [2:0] \i_mod_iq/en_gen_map/cpt ;
  wire   [4:0] \i_iq_demod/demod/QC ;
  wire   [4:0] \i_iq_demod/demod/IC ;
  wire   [4:0] \i_iq_demod/demod/QS ;
  wire   [4:0] \i_iq_demod/demod/IS ;
  wire   [17:0] \i_iq_demod/filtre_I/mult2 ;
  wire   [17:0] \i_iq_demod/filtre_I/mult1 ;
  wire   [2:0] \i_iq_demod/filtre_I/next_state ;
  wire   [17:0] \i_iq_demod/filtre_I/n_temp ;
  wire   [15:0] \i_iq_demod/filtre_I/tot ;
  wire   [17:0] \i_iq_demod/filtre_I/temp ;
  wire   [31:0] \i_iq_demod/filtre_I/current_state ;
  wire   [2:0] \i_iq_demod/filtre_I/shift_count ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg10 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg11 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg12 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg13 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg14 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg15 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg16 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg17 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg18 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg19 ;
  wire   [2:0] \i_iq_demod/filtre_I/sel ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg9 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg8 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg7 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg6 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg5 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg4 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg3 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg2 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg1 ;
  wire   [4:0] \i_iq_demod/filtre_I/shift_reg0 ;
  wire   [8:0] \i_iq_demod/filtre_I/out_factor2_req ;
  wire   [8:0] \i_iq_demod/filtre_I/out_factor1_req ;
  wire   [4:0] \i_iq_demod/filtre_I/data_2_2_req ;
  wire   [4:0] \i_iq_demod/filtre_I/data_1_2_req ;
  wire   [4:0] \i_iq_demod/filtre_I/data_2_1_req ;
  wire   [4:0] \i_iq_demod/filtre_I/data_1_1_req ;
  wire   [8:0] \i_iq_demod/filtre_I/out_factor2 ;
  wire   [8:0] \i_iq_demod/filtre_I/out_factor1 ;
  wire   [4:0] \i_iq_demod/filtre_I/data_2_2 ;
  wire   [4:0] \i_iq_demod/filtre_I/data_1_2 ;
  wire   [4:0] \i_iq_demod/filtre_I/data_2_1 ;
  wire   [4:0] \i_iq_demod/filtre_I/data_1_1 ;
  wire   [2:0] \i_iq_demod/gen_sin/next_state ;
  wire   [2:0] \i_iq_demod/gen_sin/counter ;
  wire   [31:0] \i_iq_demod/gen_sin/current_state ;
  wire   [5:0] \i_cdr/i_bit_recovery/phase_r ;
  wire   [5:0] \i_cdr/i_bit_recovery/phase_q ;
  wire   [1:0] \i_cdr/i_bit_recovery/next_state ;
  wire   [31:0] \i_cdr/i_bit_recovery/curr_state ;
  wire   [4:0] \i_cdr/i_cdr/count ;
  wire   [1:0] \i_cdr/i_cdr/next_state ;
  wire   [1:0] \i_iq_demod/demod/validation/next_state_valid ;
  wire   [31:0] \i_iq_demod/demod/validation/current_state_valid ;
  wire   [8:0] \i_iq_demod/filtre_I/mult1_multiplier/S_pipe ;
  wire   [8:0] \i_iq_demod/filtre_I/mult1_multiplier/A_pipe ;
  wire   [17:0] \i_iq_demod/filtre_Q/mult2 ;
  wire   [17:0] \i_iq_demod/filtre_Q/mult1 ;
  wire   [2:0] \i_iq_demod/filtre_Q/next_state ;
  wire   [17:0] \i_iq_demod/filtre_Q/n_temp ;
  wire   [15:0] \i_iq_demod/filtre_Q/tot ;
  wire   [17:0] \i_iq_demod/filtre_Q/temp ;
  wire   [31:0] \i_iq_demod/filtre_Q/current_state ;
  wire   [2:0] \i_iq_demod/filtre_Q/shift_count ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg10 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg11 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg12 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg13 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg14 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg15 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg16 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg17 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg18 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg19 ;
  wire   [2:0] \i_iq_demod/filtre_Q/sel ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg9 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg8 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg7 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg6 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg5 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg4 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg3 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg2 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg1 ;
  wire   [4:0] \i_iq_demod/filtre_Q/shift_reg0 ;
  wire   [8:0] \i_iq_demod/filtre_Q/out_factor2_req ;
  wire   [8:0] \i_iq_demod/filtre_Q/out_factor1_req ;
  wire   [4:0] \i_iq_demod/filtre_Q/data_2_2_req ;
  wire   [4:0] \i_iq_demod/filtre_Q/data_1_2_req ;
  wire   [4:0] \i_iq_demod/filtre_Q/data_2_1_req ;
  wire   [4:0] \i_iq_demod/filtre_Q/data_1_1_req ;
  wire   [8:0] \i_iq_demod/filtre_Q/out_factor2 ;
  wire   [8:0] \i_iq_demod/filtre_Q/out_factor1 ;
  wire   [4:0] \i_iq_demod/filtre_Q/data_2_2 ;
  wire   [4:0] \i_iq_demod/filtre_Q/data_1_2 ;
  wire   [4:0] \i_iq_demod/filtre_Q/data_2_1 ;
  wire   [4:0] \i_iq_demod/filtre_Q/data_1_1 ;
  wire   [8:0] \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe ;
  wire   [8:0] \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe ;
  wire   [8:0] \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe ;
  wire   [8:0] \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe ;
  wire   [8:0] \i_iq_demod/filtre_I/mult2_multiplier/S_pipe ;
  wire   [8:0] \i_iq_demod/filtre_I/mult2_multiplier/A_pipe ;
  wire   [4:2] \i_cdr/i_cdr/add_119/carry ;
  wire   [5:1] \i_cordic/S1/add_50/carry ;
  wire   [5:0] \i_cordic/S1/sub_50/B_not ;
  wire   [6:0] \i_cordic/S1/sub_50/carry ;
  wire   [5:0] \i_cordic/S1/sub_53/B_not ;
  wire   [6:0] \i_cordic/S1/sub_53/carry ;
  wire   [5:1] \i_cordic/S1/add_53/carry ;
  wire   [5:1] \i_cordic/S0/r64/carry ;
  wire   [5:0] \i_cordic/S0/sub_50/B_not ;
  wire   [6:0] \i_cordic/S0/sub_50/carry ;
  wire   [6:0] \i_cordic/S0/sub_53/carry ;
  wire   [5:0] \i_iq_demod/demod/r69/carry ;
  wire   [5:0] \i_iq_demod/demod/r70/carry ;
  wire   [4:0] \i_iq_demod/demod/dp_cluster_0/sub_88/B_not ;
  wire   [5:0] \i_iq_demod/demod/dp_cluster_0/sub_88/carry ;
  wire   [4:0] \i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not ;
  wire   [5:0] \i_iq_demod/demod/dp_cluster_0/sub_mult_88/carry ;
  wire   [4:1] \i_iq_demod/demod/dp_cluster_1/add_87/carry ;
  wire   [4:0] \i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not ;
  wire   [5:0] \i_iq_demod/demod/dp_cluster_1/sub_mult_87/carry ;
  wire   [7:2] \i_fifo_rx/add_90/carry ;
  wire   [6:2] \i_fifo_rx/add_106/carry ;
  wire   [6:2] \i_fifo_rx/add_139/carry ;
  wire   [5:0] \i_cordic/sub_170/carry ;
  wire   [5:0] \i_cordic/sub_173/carry ;
  wire   [4:2] \i_fifo_tx/r80/carry ;
  wire   [6:2] \i_fifo_tx/add_100/carry ;
  wire   [6:2] \i_fifo_tx/add_180/carry ;

  OAI210 U3 ( .A(N10), .B(n191), .C(n3), .Q(mux_o[9]) );
  AOI220 U4 ( .A(mod_iq_valid_o), .B(n4), .C(demod_iq_ibb_o[2]), .D(n5), .Q(n3) );
  NAND20 U5 ( .A(n6), .B(n7), .Q(mux_o[8]) );
  AOI220 U6 ( .A(fifo_rx_pslv_err_o), .B(fifo_rx_psel_i), .C(
        fifo_tx_pslv_err_o), .D(n8), .Q(n7) );
  CLKIN0 U7 ( .A(n9), .Q(n8) );
  AOI220 U8 ( .A(demod_iq_ibb_o[1]), .B(n5), .C(cdr_valid_o), .D(N13), .Q(n6)
         );
  OAI210 U9 ( .A(n191), .B(N12), .C(n11), .Q(mux_o[7]) );
  AOI220 U10 ( .A(fifo_rx_prdata_o[7]), .B(n12), .C(demod_iq_ibb_o[0]), .D(n5), 
        .Q(n11) );
  CLKIN0 U11 ( .A(n13), .Q(mux_o[6]) );
  AOI220 U12 ( .A(n12), .B(fifo_rx_prdata_o[6]), .C(n14), .D(cordic_valid_o), 
        .Q(n13) );
  CLKIN0 U13 ( .A(n15), .Q(mux_o[5]) );
  AOI220 U14 ( .A(n12), .B(fifo_rx_prdata_o[5]), .C(n14), .D(cordic_phase_o[5]), .Q(n15) );
  CLKIN0 U15 ( .A(n16), .Q(mux_o[4]) );
  AOI220 U16 ( .A(n12), .B(fifo_rx_prdata_o[4]), .C(n14), .D(cordic_phase_o[4]), .Q(n16) );
  CLKIN0 U17 ( .A(n17), .Q(mux_o[3]) );
  AOI220 U18 ( .A(n12), .B(fifo_rx_prdata_o[3]), .C(n14), .D(cordic_phase_o[3]), .Q(n17) );
  CLKIN0 U19 ( .A(n18), .Q(mux_o[2]) );
  AOI220 U20 ( .A(n12), .B(fifo_rx_prdata_o[2]), .C(n14), .D(cordic_phase_o[2]), .Q(n18) );
  CLKIN0 U21 ( .A(n19), .Q(mux_o[1]) );
  AOI220 U22 ( .A(n12), .B(fifo_rx_prdata_o[1]), .C(n14), .D(cordic_phase_o[1]), .Q(n19) );
  CLKIN0 U23 ( .A(n20), .Q(mux_o[17]) );
  AOI220 U24 ( .A(n5), .B(demod_iq_valid_o), .C(n4), .D(mod_iq_qbb_o[3]), .Q(
        n20) );
  CLKIN0 U25 ( .A(n21), .Q(mux_o[16]) );
  AOI220 U26 ( .A(n5), .B(demod_iq_qbb_o[4]), .C(n4), .D(mod_iq_qbb_o[2]), .Q(
        n21) );
  CLKIN0 U27 ( .A(n22), .Q(mux_o[15]) );
  AOI220 U28 ( .A(n5), .B(demod_iq_qbb_o[3]), .C(n4), .D(mod_iq_qbb_o[1]), .Q(
        n22) );
  CLKIN0 U29 ( .A(n23), .Q(mux_o[14]) );
  AOI220 U30 ( .A(n5), .B(demod_iq_qbb_o[2]), .C(n4), .D(mod_iq_qbb_o[0]), .Q(
        n23) );
  OAI210 U31 ( .A(N10), .B(n182), .C(n25), .Q(mux_o[13]) );
  AOI220 U32 ( .A(mod_iq_ibb_o[3]), .B(n4), .C(demod_iq_qbb_o[1]), .D(n5), .Q(
        n25) );
  OAI210 U33 ( .A(N10), .B(n286), .C(n27), .Q(mux_o[12]) );
  AOI220 U34 ( .A(mod_iq_ibb_o[2]), .B(n4), .C(demod_iq_qbb_o[0]), .D(n5), .Q(
        n27) );
  NAND20 U35 ( .A(n28), .B(n29), .Q(mux_o[11]) );
  NAND20 U36 ( .A(fifo_tx_mem_state_o), .B(N11), .Q(n29) );
  AOI220 U37 ( .A(mod_iq_ibb_o[1]), .B(n4), .C(demod_iq_ibb_o[4]), .D(n5), .Q(
        n28) );
  OAI210 U38 ( .A(N10), .B(n186), .C(n31), .Q(mux_o[10]) );
  AOI220 U39 ( .A(mod_iq_ibb_o[0]), .B(n4), .C(demod_iq_ibb_o[3]), .D(n5), .Q(
        n31) );
  CLKIN0 U41 ( .A(n33), .Q(mux_o[0]) );
  AOI220 U42 ( .A(n12), .B(fifo_rx_prdata_o[0]), .C(n14), .D(cordic_phase_o[0]), .Q(n33) );
  OAI220 U43 ( .A(N12), .B(n34), .C(n35), .D(n182), .Q(mod_iq_enable_i) );
  OAI220 U45 ( .A(N12), .B(n36), .C(n35), .D(n286), .Q(mod_iq_data_i) );
  NOR20 U47 ( .A(n12), .B(n5), .Q(n35) );
  NOR20 U48 ( .A(n9), .B(n37), .Q(fifo_tx_pwrite_i) );
  NAND20 U50 ( .A(n12), .B(mux_i[10]), .Q(n38) );
  NAND20 U52 ( .A(n12), .B(mux_i[9]), .Q(n39) );
  NAND20 U54 ( .A(n12), .B(mux_i[8]), .Q(n40) );
  NAND20 U56 ( .A(n12), .B(mux_i[7]), .Q(n41) );
  NAND20 U58 ( .A(n12), .B(mux_i[6]), .Q(n42) );
  NAND20 U60 ( .A(n12), .B(mux_i[5]), .Q(n43) );
  NAND20 U62 ( .A(n12), .B(mux_i[4]), .Q(n44) );
  NAND20 U64 ( .A(n12), .B(mux_i[3]), .Q(n45) );
  NOR20 U65 ( .A(n9), .B(n46), .Q(fifo_tx_pen_i) );
  NAND20 U66 ( .A(n48), .B(n12), .Q(n9) );
  OAI220 U67 ( .A(N10), .B(n34), .C(n47), .D(n186), .Q(fifo_rx_valid_i) );
  CLKIN0 U70 ( .A(mux_i[2]), .Q(n37) );
  CLKIN0 U72 ( .A(mux_i[1]), .Q(n46) );
  NOR20 U75 ( .A(n14), .B(n49), .Q(n47) );
  CLKIN0 U76 ( .A(n48), .Q(fifo_rx_psel_i) );
  NAND20 U77 ( .A(mux_i[0]), .B(n12), .Q(n48) );
  NOR20 U80 ( .A(n52), .B(n51), .Q(demod_iq_qif_i[4]) );
  CLKIN0 U81 ( .A(mux_i[20]), .Q(n52) );
  NOR20 U82 ( .A(n51), .B(n34), .Q(demod_iq_qif_i[3]) );
  CLKIN0 U83 ( .A(mux_i[19]), .Q(n34) );
  NOR20 U84 ( .A(n51), .B(n36), .Q(demod_iq_qif_i[2]) );
  CLKIN0 U85 ( .A(mux_i[18]), .Q(n36) );
  NOR20 U86 ( .A(n51), .B(n53), .Q(demod_iq_qif_i[1]) );
  NOR20 U87 ( .A(n51), .B(n54), .Q(\i_iq_demod/demod/N41 ) );
  NOR20 U88 ( .A(n51), .B(n55), .Q(demod_iq_iif_i[4]) );
  NOR20 U89 ( .A(n51), .B(n56), .Q(demod_iq_iif_i[3]) );
  NOR20 U90 ( .A(n51), .B(n57), .Q(demod_iq_iif_i[2]) );
  NOR20 U91 ( .A(n51), .B(n58), .Q(demod_iq_iif_i[1]) );
  NOR20 U92 ( .A(n51), .B(n59), .Q(\i_iq_demod/demod/N36 ) );
  CLKIN0 U93 ( .A(n60), .Q(cordic_valid_i) );
  AOI220 U94 ( .A(n12), .B(demod_iq_valid_o), .C(n14), .D(mux_i[10]), .Q(n60)
         );
  CLKIN0 U95 ( .A(n61), .Q(cordic_qbb_i[4]) );
  AOI220 U96 ( .A(n12), .B(demod_iq_qbb_o[4]), .C(n14), .D(mux_i[9]), .Q(n61)
         );
  CLKIN0 U97 ( .A(n62), .Q(cordic_qbb_i[3]) );
  AOI220 U98 ( .A(n12), .B(demod_iq_qbb_o[3]), .C(n14), .D(mux_i[8]), .Q(n62)
         );
  CLKIN0 U99 ( .A(n63), .Q(cordic_qbb_i[2]) );
  AOI220 U100 ( .A(n12), .B(demod_iq_qbb_o[2]), .C(n14), .D(mux_i[7]), .Q(n63)
         );
  CLKIN0 U101 ( .A(n64), .Q(cordic_qbb_i[1]) );
  AOI220 U102 ( .A(n12), .B(demod_iq_qbb_o[1]), .C(n14), .D(mux_i[6]), .Q(n64)
         );
  CLKIN0 U103 ( .A(n65), .Q(cordic_qbb_i[0]) );
  AOI220 U104 ( .A(n12), .B(demod_iq_qbb_o[0]), .C(n14), .D(mux_i[5]), .Q(n65)
         );
  CLKIN0 U105 ( .A(n66), .Q(cordic_ibb_i[4]) );
  AOI220 U106 ( .A(n12), .B(demod_iq_ibb_o[4]), .C(n14), .D(mux_i[4]), .Q(n66)
         );
  CLKIN0 U107 ( .A(n67), .Q(cordic_ibb_i[3]) );
  AOI220 U108 ( .A(n12), .B(demod_iq_ibb_o[3]), .C(n14), .D(mux_i[3]), .Q(n67)
         );
  CLKIN0 U109 ( .A(n68), .Q(cordic_ibb_i[2]) );
  AOI220 U110 ( .A(n12), .B(demod_iq_ibb_o[2]), .C(n14), .D(mux_i[2]), .Q(n68)
         );
  CLKIN0 U111 ( .A(n69), .Q(cordic_ibb_i[1]) );
  AOI220 U112 ( .A(n12), .B(demod_iq_ibb_o[1]), .C(n14), .D(mux_i[1]), .Q(n69)
         );
  CLKIN0 U113 ( .A(n70), .Q(cordic_ibb_i[0]) );
  AOI220 U114 ( .A(n12), .B(demod_iq_ibb_o[0]), .C(n14), .D(mux_i[0]), .Q(n70)
         );
  OAI220 U119 ( .A(n51), .B(n251), .C(n73), .D(n53), .Q(cdr_valid_i) );
  CLKIN0 U120 ( .A(mux_i[17]), .Q(n53) );
  OAI220 U122 ( .A(n51), .B(n258), .C(n73), .D(n54), .Q(cdr_phase_i[5]) );
  CLKIN0 U123 ( .A(mux_i[16]), .Q(n54) );
  OAI220 U125 ( .A(n51), .B(n257), .C(n73), .D(n55), .Q(cdr_phase_i[4]) );
  CLKIN0 U126 ( .A(mux_i[15]), .Q(n55) );
  OAI220 U128 ( .A(n51), .B(n256), .C(n73), .D(n56), .Q(cdr_phase_i[3]) );
  CLKIN0 U129 ( .A(mux_i[14]), .Q(n56) );
  OAI220 U131 ( .A(n51), .B(n255), .C(n73), .D(n57), .Q(cdr_phase_i[2]) );
  CLKIN0 U132 ( .A(mux_i[13]), .Q(n57) );
  OAI220 U134 ( .A(n51), .B(n254), .C(n73), .D(n58), .Q(cdr_phase_i[1]) );
  CLKIN0 U135 ( .A(mux_i[12]), .Q(n58) );
  OAI220 U137 ( .A(n51), .B(n253), .C(n73), .D(n59), .Q(cdr_phase_i[0]) );
  CLKIN0 U138 ( .A(mux_i[11]), .Q(n59) );
  NAND20 U143 ( .A(sel_i[1]), .B(sel_i[0]), .Q(n71) );
  NAND20 U145 ( .A(n80), .B(n81), .Q(n32) );
  CLKIN0 U147 ( .A(sel_i[0]), .Q(n80) );
  CLKIN0 U149 ( .A(sel_i[1]), .Q(n81) );
  NOR30 \i_fifo_tx/U205  ( .A(\i_fifo_tx/counter_clock [0]), .B(
        \i_fifo_tx/counter_clock [2]), .C(\i_fifo_tx/counter_clock [1]), .Q(
        \i_fifo_tx/n203 ) );
  NOR20 \i_fifo_tx/U201  ( .A(\i_fifo_tx/n81 ), .B(
        \i_fifo_tx/counter_clock [0]), .Q(\i_fifo_tx/N187 ) );
  CLKIN0 \i_fifo_tx/U200  ( .A(\i_fifo_tx/N149 ), .Q(\i_fifo_tx/n201 ) );
  NOR20 \i_fifo_tx/U199  ( .A(\i_fifo_tx/n81 ), .B(\i_fifo_tx/n201 ), .Q(
        \i_fifo_tx/N188 ) );
  CLKIN0 \i_fifo_tx/U198  ( .A(\i_fifo_tx/N150 ), .Q(\i_fifo_tx/n200 ) );
  NOR20 \i_fifo_tx/U197  ( .A(\i_fifo_tx/n81 ), .B(\i_fifo_tx/n200 ), .Q(
        \i_fifo_tx/N189 ) );
  CLKIN0 \i_fifo_tx/U196  ( .A(\i_fifo_tx/N151 ), .Q(\i_fifo_tx/n199 ) );
  NOR20 \i_fifo_tx/U195  ( .A(\i_fifo_tx/n81 ), .B(\i_fifo_tx/n199 ), .Q(
        \i_fifo_tx/N190 ) );
  NOR20 \i_fifo_tx/U193  ( .A(\i_fifo_tx/n81 ), .B(n245), .Q(\i_fifo_tx/N191 )
         );
  XNR20 \i_fifo_tx/U190  ( .A(\i_fifo_tx/n183 ), .B(\i_fifo_tx/n188 ), .Q(
        \i_fifo_tx/n186 ) );
  NAND20 \i_fifo_tx/U189  ( .A(\i_fifo_tx/n186 ), .B(\i_fifo_tx/N40 ), .Q(
        fifo_tx_mem_state_o) );
  NAND30 \i_fifo_tx/U188  ( .A(\i_fifo_tx/N37 ), .B(\i_fifo_tx/N36 ), .C(
        \i_fifo_tx/N38 ), .Q(\i_fifo_tx/n189 ) );
  NAND20 \i_fifo_tx/U187  ( .A(\i_fifo_tx/state_rd ), .B(\i_fifo_tx/n189 ), 
        .Q(\i_fifo_tx/n194 ) );
  NAND20 \i_fifo_tx/U186  ( .A(\i_fifo_tx/n81 ), .B(\i_fifo_tx/n195 ), .Q(
        \i_fifo_tx/n196 ) );
  OAI220 \i_fifo_tx/U185  ( .A(\i_fifo_tx/n81 ), .B(\i_fifo_tx/n195 ), .C(
        \i_fifo_tx/n194 ), .D(\i_fifo_tx/n196 ), .Q(\i_fifo_tx/n207 ) );
  CLKIN0 \i_fifo_tx/U184  ( .A(\i_fifo_tx/n194 ), .Q(\i_fifo_tx/n85 ) );
  OAI210 \i_fifo_tx/U183  ( .A(\i_fifo_tx/N36 ), .B(\i_fifo_tx/n194 ), .C(
        \i_fifo_tx/n81 ), .Q(\i_fifo_tx/n86 ) );
  OAI210 \i_fifo_tx/U182  ( .A(\i_fifo_tx/n85 ), .B(\i_fifo_tx/n86 ), .C(
        \i_fifo_tx/N38 ), .Q(\i_fifo_tx/n192 ) );
  NAND40 \i_fifo_tx/U181  ( .A(\i_fifo_tx/n85 ), .B(\i_fifo_tx/N37 ), .C(
        \i_fifo_tx/N36 ), .D(\i_fifo_tx/n81 ), .Q(\i_fifo_tx/n193 ) );
  NAND20 \i_fifo_tx/U180  ( .A(\i_fifo_tx/n192 ), .B(\i_fifo_tx/n193 ), .Q(
        \i_fifo_tx/n206 ) );
  CLKIN0 \i_fifo_tx/U178  ( .A(\i_fifo_tx/N40 ), .Q(\i_fifo_tx/n185 ) );
  NOR20 \i_fifo_tx/U177  ( .A(\i_fifo_tx/n185 ), .B(\i_fifo_tx/n186 ), .Q(
        fifo_tx_pslv_err_o) );
  NAND20 \i_fifo_tx/U170  ( .A(\i_fifo_tx/n179 ), .B(\i_fifo_tx/n169 ), .Q(
        \i_fifo_tx/n151 ) );
  NAND20 \i_fifo_tx/U168  ( .A(\i_fifo_tx/n179 ), .B(\i_fifo_tx/n168 ), .Q(
        \i_fifo_tx/n150 ) );
  NAND20 \i_fifo_tx/U166  ( .A(\i_fifo_tx/n179 ), .B(\i_fifo_tx/n167 ), .Q(
        \i_fifo_tx/n149 ) );
  NAND20 \i_fifo_tx/U164  ( .A(\i_fifo_tx/n179 ), .B(\i_fifo_tx/n166 ), .Q(
        \i_fifo_tx/n148 ) );
  NAND20 \i_fifo_tx/U162  ( .A(\i_fifo_tx/n179 ), .B(\i_fifo_tx/n165 ), .Q(
        \i_fifo_tx/n147 ) );
  NAND20 \i_fifo_tx/U160  ( .A(\i_fifo_tx/n179 ), .B(\i_fifo_tx/n164 ), .Q(
        \i_fifo_tx/n146 ) );
  NAND20 \i_fifo_tx/U158  ( .A(\i_fifo_tx/n179 ), .B(\i_fifo_tx/n163 ), .Q(
        \i_fifo_tx/n145 ) );
  NAND20 \i_fifo_tx/U156  ( .A(\i_fifo_tx/n179 ), .B(\i_fifo_tx/n162 ), .Q(
        \i_fifo_tx/n144 ) );
  NAND20 \i_fifo_tx/U154  ( .A(\i_fifo_tx/n178 ), .B(\i_fifo_tx/n169 ), .Q(
        \i_fifo_tx/n143 ) );
  NAND20 \i_fifo_tx/U153  ( .A(\i_fifo_tx/n178 ), .B(\i_fifo_tx/n168 ), .Q(
        \i_fifo_tx/n142 ) );
  NAND20 \i_fifo_tx/U152  ( .A(\i_fifo_tx/n178 ), .B(\i_fifo_tx/n167 ), .Q(
        \i_fifo_tx/n141 ) );
  NAND20 \i_fifo_tx/U151  ( .A(\i_fifo_tx/n178 ), .B(\i_fifo_tx/n166 ), .Q(
        \i_fifo_tx/n140 ) );
  NAND20 \i_fifo_tx/U150  ( .A(\i_fifo_tx/n178 ), .B(\i_fifo_tx/n165 ), .Q(
        \i_fifo_tx/n139 ) );
  NAND20 \i_fifo_tx/U149  ( .A(\i_fifo_tx/n178 ), .B(\i_fifo_tx/n164 ), .Q(
        \i_fifo_tx/n138 ) );
  NAND20 \i_fifo_tx/U148  ( .A(\i_fifo_tx/n178 ), .B(\i_fifo_tx/n163 ), .Q(
        \i_fifo_tx/n137 ) );
  NAND20 \i_fifo_tx/U147  ( .A(\i_fifo_tx/n178 ), .B(\i_fifo_tx/n162 ), .Q(
        \i_fifo_tx/n136 ) );
  NAND20 \i_fifo_tx/U145  ( .A(\i_fifo_tx/n177 ), .B(\i_fifo_tx/n169 ), .Q(
        \i_fifo_tx/n135 ) );
  NAND20 \i_fifo_tx/U144  ( .A(\i_fifo_tx/n177 ), .B(\i_fifo_tx/n168 ), .Q(
        \i_fifo_tx/n134 ) );
  NAND20 \i_fifo_tx/U143  ( .A(\i_fifo_tx/n177 ), .B(\i_fifo_tx/n167 ), .Q(
        \i_fifo_tx/n133 ) );
  NAND20 \i_fifo_tx/U142  ( .A(\i_fifo_tx/n177 ), .B(\i_fifo_tx/n166 ), .Q(
        \i_fifo_tx/n132 ) );
  NAND20 \i_fifo_tx/U141  ( .A(\i_fifo_tx/n177 ), .B(\i_fifo_tx/n165 ), .Q(
        \i_fifo_tx/n131 ) );
  NAND20 \i_fifo_tx/U140  ( .A(\i_fifo_tx/n177 ), .B(\i_fifo_tx/n164 ), .Q(
        \i_fifo_tx/n130 ) );
  NAND20 \i_fifo_tx/U139  ( .A(\i_fifo_tx/n177 ), .B(\i_fifo_tx/n163 ), .Q(
        \i_fifo_tx/n129 ) );
  NAND20 \i_fifo_tx/U138  ( .A(\i_fifo_tx/n177 ), .B(\i_fifo_tx/n162 ), .Q(
        \i_fifo_tx/n128 ) );
  NAND20 \i_fifo_tx/U136  ( .A(\i_fifo_tx/n176 ), .B(\i_fifo_tx/n169 ), .Q(
        \i_fifo_tx/n127 ) );
  NAND20 \i_fifo_tx/U135  ( .A(\i_fifo_tx/n176 ), .B(\i_fifo_tx/n168 ), .Q(
        \i_fifo_tx/n126 ) );
  NAND20 \i_fifo_tx/U134  ( .A(\i_fifo_tx/n176 ), .B(\i_fifo_tx/n167 ), .Q(
        \i_fifo_tx/n125 ) );
  NAND20 \i_fifo_tx/U133  ( .A(\i_fifo_tx/n176 ), .B(\i_fifo_tx/n166 ), .Q(
        \i_fifo_tx/n124 ) );
  NAND20 \i_fifo_tx/U132  ( .A(\i_fifo_tx/n176 ), .B(\i_fifo_tx/n165 ), .Q(
        \i_fifo_tx/n123 ) );
  NAND20 \i_fifo_tx/U131  ( .A(\i_fifo_tx/n176 ), .B(\i_fifo_tx/n164 ), .Q(
        \i_fifo_tx/n122 ) );
  NAND20 \i_fifo_tx/U130  ( .A(\i_fifo_tx/n176 ), .B(\i_fifo_tx/n163 ), .Q(
        \i_fifo_tx/n121 ) );
  NAND20 \i_fifo_tx/U129  ( .A(\i_fifo_tx/n176 ), .B(\i_fifo_tx/n162 ), .Q(
        \i_fifo_tx/n120 ) );
  NAND20 \i_fifo_tx/U127  ( .A(\i_fifo_tx/n175 ), .B(\i_fifo_tx/n169 ), .Q(
        \i_fifo_tx/n119 ) );
  NAND20 \i_fifo_tx/U126  ( .A(\i_fifo_tx/n175 ), .B(\i_fifo_tx/n168 ), .Q(
        \i_fifo_tx/n118 ) );
  NAND20 \i_fifo_tx/U125  ( .A(\i_fifo_tx/n175 ), .B(\i_fifo_tx/n167 ), .Q(
        \i_fifo_tx/n117 ) );
  NAND20 \i_fifo_tx/U124  ( .A(\i_fifo_tx/n175 ), .B(\i_fifo_tx/n166 ), .Q(
        \i_fifo_tx/n116 ) );
  NAND20 \i_fifo_tx/U123  ( .A(\i_fifo_tx/n175 ), .B(\i_fifo_tx/n165 ), .Q(
        \i_fifo_tx/n115 ) );
  NAND20 \i_fifo_tx/U122  ( .A(\i_fifo_tx/n175 ), .B(\i_fifo_tx/n164 ), .Q(
        \i_fifo_tx/n114 ) );
  NAND20 \i_fifo_tx/U121  ( .A(\i_fifo_tx/n175 ), .B(\i_fifo_tx/n163 ), .Q(
        \i_fifo_tx/n113 ) );
  NAND20 \i_fifo_tx/U120  ( .A(\i_fifo_tx/n175 ), .B(\i_fifo_tx/n162 ), .Q(
        \i_fifo_tx/n112 ) );
  NAND20 \i_fifo_tx/U118  ( .A(\i_fifo_tx/n174 ), .B(\i_fifo_tx/n169 ), .Q(
        \i_fifo_tx/n111 ) );
  NAND20 \i_fifo_tx/U117  ( .A(\i_fifo_tx/n174 ), .B(\i_fifo_tx/n168 ), .Q(
        \i_fifo_tx/n110 ) );
  NAND20 \i_fifo_tx/U116  ( .A(\i_fifo_tx/n174 ), .B(\i_fifo_tx/n167 ), .Q(
        \i_fifo_tx/n109 ) );
  NAND20 \i_fifo_tx/U115  ( .A(\i_fifo_tx/n174 ), .B(\i_fifo_tx/n166 ), .Q(
        \i_fifo_tx/n108 ) );
  NAND20 \i_fifo_tx/U114  ( .A(\i_fifo_tx/n174 ), .B(\i_fifo_tx/n165 ), .Q(
        \i_fifo_tx/n107 ) );
  NAND20 \i_fifo_tx/U113  ( .A(\i_fifo_tx/n174 ), .B(\i_fifo_tx/n164 ), .Q(
        \i_fifo_tx/n106 ) );
  NAND20 \i_fifo_tx/U112  ( .A(\i_fifo_tx/n174 ), .B(\i_fifo_tx/n163 ), .Q(
        \i_fifo_tx/n105 ) );
  NAND20 \i_fifo_tx/U111  ( .A(\i_fifo_tx/n174 ), .B(\i_fifo_tx/n162 ), .Q(
        \i_fifo_tx/n104 ) );
  NAND20 \i_fifo_tx/U109  ( .A(\i_fifo_tx/n173 ), .B(\i_fifo_tx/n169 ), .Q(
        \i_fifo_tx/n103 ) );
  NAND20 \i_fifo_tx/U108  ( .A(\i_fifo_tx/n173 ), .B(\i_fifo_tx/n168 ), .Q(
        \i_fifo_tx/n102 ) );
  NAND20 \i_fifo_tx/U107  ( .A(\i_fifo_tx/n173 ), .B(\i_fifo_tx/n167 ), .Q(
        \i_fifo_tx/n101 ) );
  NAND20 \i_fifo_tx/U106  ( .A(\i_fifo_tx/n173 ), .B(\i_fifo_tx/n166 ), .Q(
        \i_fifo_tx/n100 ) );
  NAND20 \i_fifo_tx/U105  ( .A(\i_fifo_tx/n173 ), .B(\i_fifo_tx/n165 ), .Q(
        \i_fifo_tx/n99 ) );
  NAND20 \i_fifo_tx/U104  ( .A(\i_fifo_tx/n173 ), .B(\i_fifo_tx/n164 ), .Q(
        \i_fifo_tx/n98 ) );
  NAND20 \i_fifo_tx/U103  ( .A(\i_fifo_tx/n173 ), .B(\i_fifo_tx/n163 ), .Q(
        \i_fifo_tx/n97 ) );
  NAND20 \i_fifo_tx/U102  ( .A(\i_fifo_tx/n173 ), .B(\i_fifo_tx/n162 ), .Q(
        \i_fifo_tx/n96 ) );
  NAND20 \i_fifo_tx/U100  ( .A(\i_fifo_tx/n169 ), .B(\i_fifo_tx/n161 ), .Q(
        \i_fifo_tx/n95 ) );
  NAND20 \i_fifo_tx/U99  ( .A(\i_fifo_tx/n168 ), .B(\i_fifo_tx/n161 ), .Q(
        \i_fifo_tx/n94 ) );
  NAND20 \i_fifo_tx/U98  ( .A(\i_fifo_tx/n167 ), .B(\i_fifo_tx/n161 ), .Q(
        \i_fifo_tx/n93 ) );
  NAND20 \i_fifo_tx/U97  ( .A(\i_fifo_tx/n166 ), .B(\i_fifo_tx/n161 ), .Q(
        \i_fifo_tx/n92 ) );
  NAND20 \i_fifo_tx/U96  ( .A(\i_fifo_tx/n165 ), .B(\i_fifo_tx/n161 ), .Q(
        \i_fifo_tx/n91 ) );
  NAND20 \i_fifo_tx/U95  ( .A(\i_fifo_tx/n164 ), .B(\i_fifo_tx/n161 ), .Q(
        \i_fifo_tx/n90 ) );
  NAND20 \i_fifo_tx/U94  ( .A(\i_fifo_tx/n163 ), .B(\i_fifo_tx/n161 ), .Q(
        \i_fifo_tx/n89 ) );
  NAND20 \i_fifo_tx/U93  ( .A(\i_fifo_tx/n161 ), .B(\i_fifo_tx/n162 ), .Q(
        \i_fifo_tx/n88 ) );
  CLKIN0 \i_fifo_tx/U85  ( .A(\i_fifo_tx/n86 ), .Q(\i_fifo_tx/n82 ) );
  NAND40 \i_fifo_tx/U84  ( .A(\i_fifo_tx/n85 ), .B(\i_fifo_tx/N36 ), .C(
        \i_fifo_tx/n81 ), .D(\i_fifo_tx/n83 ), .Q(\i_fifo_tx/n84 ) );
  OAI210 \i_fifo_tx/U83  ( .A(\i_fifo_tx/n82 ), .B(\i_fifo_tx/n83 ), .C(
        \i_fifo_tx/n84 ), .Q(\i_fifo_tx/n205 ) );
  NAND30 \i_fifo_tx/U81  ( .A(\i_fifo_tx/counter_clock [0]), .B(
        \i_fifo_tx/state_rd ), .C(\i_fifo_tx/counter_clock [2]), .Q(
        \i_fifo_tx/n79 ) );
  NOR40 \i_fifo_tx/U80  ( .A(\i_fifo_tx/n79 ), .B(\i_fifo_tx/n80 ), .C(
        \i_fifo_tx/counter_clock [4]), .D(\i_fifo_tx/counter_clock [1]), .Q(
        \i_fifo_tx/n78 ) );
  INV2 \i_fifo_tx/U75  ( .A(\i_fifo_tx/n127 ), .Q(\i_fifo_tx/n74 ) );
  INV2 \i_fifo_tx/U73  ( .A(\i_fifo_tx/n88 ), .Q(\i_fifo_tx/n72 ) );
  INV2 \i_fifo_tx/U72  ( .A(\i_fifo_tx/n89 ), .Q(\i_fifo_tx/n71 ) );
  INV2 \i_fifo_tx/U71  ( .A(\i_fifo_tx/n90 ), .Q(\i_fifo_tx/n70 ) );
  INV2 \i_fifo_tx/U70  ( .A(\i_fifo_tx/n91 ), .Q(\i_fifo_tx/n69 ) );
  INV2 \i_fifo_tx/U69  ( .A(\i_fifo_tx/n92 ), .Q(\i_fifo_tx/n68 ) );
  INV2 \i_fifo_tx/U68  ( .A(\i_fifo_tx/n93 ), .Q(\i_fifo_tx/n67 ) );
  INV2 \i_fifo_tx/U67  ( .A(\i_fifo_tx/n94 ), .Q(\i_fifo_tx/n66 ) );
  INV2 \i_fifo_tx/U66  ( .A(\i_fifo_tx/n95 ), .Q(\i_fifo_tx/n65 ) );
  INV2 \i_fifo_tx/U65  ( .A(\i_fifo_tx/n96 ), .Q(\i_fifo_tx/n64 ) );
  INV2 \i_fifo_tx/U64  ( .A(\i_fifo_tx/n97 ), .Q(\i_fifo_tx/n63 ) );
  INV2 \i_fifo_tx/U63  ( .A(\i_fifo_tx/n98 ), .Q(\i_fifo_tx/n62 ) );
  INV2 \i_fifo_tx/U62  ( .A(\i_fifo_tx/n99 ), .Q(\i_fifo_tx/n61 ) );
  INV2 \i_fifo_tx/U61  ( .A(\i_fifo_tx/n100 ), .Q(\i_fifo_tx/n60 ) );
  INV2 \i_fifo_tx/U60  ( .A(\i_fifo_tx/n101 ), .Q(\i_fifo_tx/n59 ) );
  INV2 \i_fifo_tx/U59  ( .A(\i_fifo_tx/n102 ), .Q(\i_fifo_tx/n58 ) );
  INV2 \i_fifo_tx/U58  ( .A(\i_fifo_tx/n103 ), .Q(\i_fifo_tx/n57 ) );
  INV2 \i_fifo_tx/U57  ( .A(\i_fifo_tx/n104 ), .Q(\i_fifo_tx/n56 ) );
  INV2 \i_fifo_tx/U56  ( .A(\i_fifo_tx/n105 ), .Q(\i_fifo_tx/n55 ) );
  INV2 \i_fifo_tx/U55  ( .A(\i_fifo_tx/n106 ), .Q(\i_fifo_tx/n54 ) );
  INV2 \i_fifo_tx/U54  ( .A(\i_fifo_tx/n107 ), .Q(\i_fifo_tx/n53 ) );
  INV2 \i_fifo_tx/U53  ( .A(\i_fifo_tx/n108 ), .Q(\i_fifo_tx/n52 ) );
  INV2 \i_fifo_tx/U52  ( .A(\i_fifo_tx/n109 ), .Q(\i_fifo_tx/n51 ) );
  INV2 \i_fifo_tx/U51  ( .A(\i_fifo_tx/n110 ), .Q(\i_fifo_tx/n50 ) );
  INV2 \i_fifo_tx/U50  ( .A(\i_fifo_tx/n111 ), .Q(\i_fifo_tx/n49 ) );
  INV2 \i_fifo_tx/U49  ( .A(\i_fifo_tx/n112 ), .Q(\i_fifo_tx/n48 ) );
  INV2 \i_fifo_tx/U48  ( .A(\i_fifo_tx/n113 ), .Q(\i_fifo_tx/n47 ) );
  INV2 \i_fifo_tx/U47  ( .A(\i_fifo_tx/n114 ), .Q(\i_fifo_tx/n46 ) );
  INV2 \i_fifo_tx/U46  ( .A(\i_fifo_tx/n115 ), .Q(\i_fifo_tx/n45 ) );
  INV2 \i_fifo_tx/U45  ( .A(\i_fifo_tx/n116 ), .Q(\i_fifo_tx/n44 ) );
  INV2 \i_fifo_tx/U44  ( .A(\i_fifo_tx/n117 ), .Q(\i_fifo_tx/n43 ) );
  INV2 \i_fifo_tx/U43  ( .A(\i_fifo_tx/n118 ), .Q(\i_fifo_tx/n42 ) );
  INV2 \i_fifo_tx/U42  ( .A(\i_fifo_tx/n119 ), .Q(\i_fifo_tx/n41 ) );
  INV2 \i_fifo_tx/U41  ( .A(\i_fifo_tx/n120 ), .Q(\i_fifo_tx/n40 ) );
  INV2 \i_fifo_tx/U40  ( .A(\i_fifo_tx/n121 ), .Q(\i_fifo_tx/n39 ) );
  INV2 \i_fifo_tx/U39  ( .A(\i_fifo_tx/n122 ), .Q(\i_fifo_tx/n38 ) );
  INV2 \i_fifo_tx/U38  ( .A(\i_fifo_tx/n123 ), .Q(\i_fifo_tx/n37 ) );
  INV2 \i_fifo_tx/U37  ( .A(\i_fifo_tx/n124 ), .Q(\i_fifo_tx/n36 ) );
  INV2 \i_fifo_tx/U36  ( .A(\i_fifo_tx/n125 ), .Q(\i_fifo_tx/n35 ) );
  INV2 \i_fifo_tx/U35  ( .A(\i_fifo_tx/n126 ), .Q(\i_fifo_tx/n34 ) );
  INV2 \i_fifo_tx/U34  ( .A(\i_fifo_tx/n128 ), .Q(\i_fifo_tx/n33 ) );
  INV2 \i_fifo_tx/U33  ( .A(\i_fifo_tx/n129 ), .Q(\i_fifo_tx/n32 ) );
  INV2 \i_fifo_tx/U32  ( .A(\i_fifo_tx/n130 ), .Q(\i_fifo_tx/n31 ) );
  INV2 \i_fifo_tx/U31  ( .A(\i_fifo_tx/n131 ), .Q(\i_fifo_tx/n30 ) );
  INV2 \i_fifo_tx/U30  ( .A(\i_fifo_tx/n132 ), .Q(\i_fifo_tx/n29 ) );
  INV2 \i_fifo_tx/U29  ( .A(\i_fifo_tx/n133 ), .Q(\i_fifo_tx/n28 ) );
  INV2 \i_fifo_tx/U28  ( .A(\i_fifo_tx/n134 ), .Q(\i_fifo_tx/n27 ) );
  INV2 \i_fifo_tx/U27  ( .A(\i_fifo_tx/n135 ), .Q(\i_fifo_tx/n26 ) );
  INV2 \i_fifo_tx/U26  ( .A(\i_fifo_tx/n136 ), .Q(\i_fifo_tx/n25 ) );
  INV2 \i_fifo_tx/U25  ( .A(\i_fifo_tx/n137 ), .Q(\i_fifo_tx/n24 ) );
  INV2 \i_fifo_tx/U24  ( .A(\i_fifo_tx/n138 ), .Q(\i_fifo_tx/n23 ) );
  INV2 \i_fifo_tx/U23  ( .A(\i_fifo_tx/n139 ), .Q(\i_fifo_tx/n22 ) );
  INV2 \i_fifo_tx/U22  ( .A(\i_fifo_tx/n140 ), .Q(\i_fifo_tx/n21 ) );
  INV2 \i_fifo_tx/U21  ( .A(\i_fifo_tx/n141 ), .Q(\i_fifo_tx/n20 ) );
  INV2 \i_fifo_tx/U20  ( .A(\i_fifo_tx/n142 ), .Q(\i_fifo_tx/n19 ) );
  INV2 \i_fifo_tx/U19  ( .A(\i_fifo_tx/n143 ), .Q(\i_fifo_tx/n18 ) );
  INV2 \i_fifo_tx/U18  ( .A(\i_fifo_tx/n144 ), .Q(\i_fifo_tx/n17 ) );
  INV2 \i_fifo_tx/U17  ( .A(\i_fifo_tx/n145 ), .Q(\i_fifo_tx/n16 ) );
  INV2 \i_fifo_tx/U16  ( .A(\i_fifo_tx/n146 ), .Q(\i_fifo_tx/n15 ) );
  INV2 \i_fifo_tx/U15  ( .A(\i_fifo_tx/n147 ), .Q(\i_fifo_tx/n14 ) );
  INV2 \i_fifo_tx/U14  ( .A(\i_fifo_tx/n148 ), .Q(\i_fifo_tx/n13 ) );
  INV2 \i_fifo_tx/U13  ( .A(\i_fifo_tx/n149 ), .Q(\i_fifo_tx/n12 ) );
  INV2 \i_fifo_tx/U12  ( .A(\i_fifo_tx/n150 ), .Q(\i_fifo_tx/n11 ) );
  INV2 \i_fifo_tx/U11  ( .A(\i_fifo_tx/n151 ), .Q(\i_fifo_tx/n10 ) );
  DFC1 \i_fifo_tx/IQ_rate_reg  ( .D(\i_fifo_tx/n204 ), .C(clk_i), .RN(resetn_i), .Q(fifo_tx_enable_o), .QN(n182) );
  DFC1 \i_fifo_tx/counter_clock_reg[4]  ( .D(\i_fifo_tx/N191 ), .C(clk_i), 
        .RN(resetn_i), .Q(\i_fifo_tx/counter_clock [4]) );
  DFC3 \i_fifo_tx/counter_clock_reg[3]  ( .D(\i_fifo_tx/N190 ), .C(clk_i), 
        .RN(resetn_i), .Q(\i_fifo_tx/counter_clock [3]), .QN(\i_fifo_tx/n80 )
         );
  DFC1 \i_fifo_tx/counter_clock_reg[2]  ( .D(\i_fifo_tx/N189 ), .C(clk_i), 
        .RN(resetn_i), .Q(\i_fifo_tx/counter_clock [2]) );
  DFC1 \i_fifo_tx/counter_clock_reg[1]  ( .D(\i_fifo_tx/N188 ), .C(clk_i), 
        .RN(resetn_i), .Q(\i_fifo_tx/counter_clock [1]) );
  DFC1 \i_fifo_tx/counter_clock_reg[0]  ( .D(\i_fifo_tx/N187 ), .C(clk_i), 
        .RN(resetn_i), .Q(\i_fifo_tx/counter_clock [0]) );
  DFC1 \i_fifo_tx/state_rd_reg  ( .D(\i_fifo_tx/next_state_rd ), .C(clk_i), 
        .RN(resetn_i), .Q(\i_fifo_tx/state_rd ), .QN(\i_fifo_tx/n190 ) );
  DFEC1 \i_fifo_tx/mem_reg[0][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n10 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[0][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[1][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n11 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[1][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[2][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[2][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[3][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n13 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[3][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[4][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n14 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[4][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[5][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n15 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[5][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[6][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n16 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[6][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[7][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n17 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[7][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[8][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n18 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[8][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[9][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n19 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[9][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[10][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n20 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[10][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[11][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n21 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[11][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[12][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n22 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[12][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[13][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n23 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[13][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[14][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[14][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[15][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n25 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[15][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[16][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n26 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[16][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[17][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[17][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[18][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n28 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[18][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[19][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n29 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[19][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[20][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[20][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[21][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n31 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[21][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[22][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n32 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[22][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[23][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[23][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[25][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n34 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[25][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[26][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n35 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[26][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[27][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[27][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[28][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n37 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[28][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[29][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n38 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[29][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[30][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[30][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[31][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n40 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[31][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[32][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n41 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[32][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[33][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[33][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[34][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n43 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[34][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[35][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n44 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[35][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[36][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n45 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[36][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[37][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n46 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[37][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[38][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n47 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[38][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[39][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[39][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[40][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n49 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[40][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[41][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n50 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[41][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[42][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[42][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[43][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n52 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[43][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[44][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[44][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[45][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n54 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[45][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[46][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[46][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[47][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n56 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[47][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[48][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[48][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[49][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n58 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[49][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[50][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[50][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[51][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n60 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[51][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[52][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[52][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[53][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n62 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[53][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[54][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[54][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[55][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n64 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[55][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[56][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[56][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[57][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n66 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[57][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[58][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n67 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[58][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[59][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[59][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[60][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n69 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[60][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[61][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[61][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[62][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n71 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[62][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[63][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[63][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[24][0]  ( .D(\i_fifo_tx/n3 ), .E(\i_fifo_tx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[24][0] ) );
  DFEC1 \i_fifo_tx/mem_reg[0][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n10 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[0][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[1][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n11 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[1][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[2][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[2][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[3][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n13 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[3][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[4][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n14 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[4][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[5][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n15 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[5][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[6][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n16 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[6][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[7][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n17 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[7][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[8][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n18 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[8][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[9][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n19 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[9][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[10][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n20 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[10][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[11][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n21 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[11][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[12][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n22 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[12][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[13][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n23 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[13][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[14][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[14][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[15][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n25 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[15][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[16][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n26 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[16][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[17][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[17][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[18][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n28 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[18][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[19][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n29 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[19][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[20][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[20][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[21][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n31 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[21][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[22][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n32 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[22][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[23][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[23][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[25][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n34 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[25][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[26][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n35 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[26][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[27][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[27][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[28][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n37 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[28][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[29][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n38 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[29][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[30][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[30][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[31][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n40 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[31][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[32][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n41 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[32][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[33][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[33][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[34][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n43 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[34][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[35][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n44 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[35][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[36][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n45 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[36][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[37][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n46 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[37][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[38][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n47 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[38][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[39][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[39][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[40][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n49 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[40][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[41][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n50 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[41][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[42][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[42][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[43][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n52 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[43][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[44][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[44][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[45][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n54 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[45][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[46][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[46][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[47][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n56 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[47][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[48][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[48][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[49][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n58 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[49][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[50][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[50][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[51][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n60 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[51][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[52][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[52][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[53][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n62 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[53][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[54][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[54][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[55][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n64 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[55][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[56][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[56][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[57][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n66 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[57][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[58][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n67 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[58][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[59][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[59][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[60][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n69 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[60][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[61][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[61][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[62][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n71 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[62][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[63][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[63][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[24][1]  ( .D(\i_fifo_tx/n4 ), .E(\i_fifo_tx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[24][1] ) );
  DFEC1 \i_fifo_tx/mem_reg[0][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n10 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[0][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[1][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n11 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[1][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[2][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[2][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[3][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n13 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[3][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[4][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n14 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[4][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[5][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n15 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[5][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[6][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n16 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[6][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[7][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n17 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[7][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[8][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n18 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[8][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[9][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n19 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[9][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[10][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n20 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[10][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[11][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n21 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[11][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[12][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n22 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[12][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[13][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n23 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[13][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[14][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[14][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[15][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n25 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[15][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[16][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n26 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[16][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[17][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[17][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[18][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n28 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[18][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[19][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n29 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[19][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[20][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[20][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[21][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n31 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[21][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[22][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n32 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[22][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[23][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[23][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[25][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n34 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[25][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[26][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n35 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[26][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[27][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[27][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[28][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n37 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[28][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[29][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n38 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[29][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[30][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[30][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[31][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n40 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[31][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[32][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n41 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[32][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[33][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[33][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[34][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n43 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[34][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[35][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n44 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[35][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[36][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n45 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[36][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[37][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n46 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[37][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[38][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n47 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[38][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[39][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[39][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[40][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n49 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[40][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[41][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n50 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[41][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[42][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[42][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[43][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n52 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[43][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[44][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[44][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[45][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n54 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[45][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[46][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[46][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[47][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n56 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[47][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[48][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[48][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[49][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n58 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[49][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[50][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[50][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[51][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n60 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[51][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[52][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[52][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[53][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n62 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[53][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[54][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[54][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[55][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n64 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[55][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[56][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[56][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[57][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n66 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[57][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[58][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n67 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[58][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[59][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[59][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[60][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n69 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[60][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[61][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[61][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[62][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n71 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[62][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[63][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[63][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[24][2]  ( .D(\i_fifo_tx/n5 ), .E(\i_fifo_tx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[24][2] ) );
  DFEC1 \i_fifo_tx/mem_reg[0][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n10 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[0][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[1][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n11 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[1][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[2][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[2][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[3][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n13 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[3][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[4][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n14 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[4][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[5][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n15 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[5][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[6][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n16 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[6][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[7][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n17 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[7][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[8][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n18 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[8][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[9][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n19 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[9][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[10][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n20 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[10][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[11][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n21 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[11][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[12][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n22 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[12][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[13][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n23 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[13][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[14][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[14][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[15][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n25 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[15][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[16][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n26 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[16][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[17][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[17][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[18][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n28 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[18][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[19][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n29 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[19][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[20][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[20][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[21][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n31 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[21][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[22][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n32 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[22][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[23][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[23][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[25][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n34 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[25][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[26][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n35 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[26][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[27][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[27][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[28][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n37 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[28][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[29][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n38 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[29][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[30][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[30][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[31][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n40 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[31][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[32][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n41 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[32][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[33][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[33][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[34][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n43 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[34][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[35][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n44 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[35][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[36][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n45 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[36][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[37][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n46 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[37][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[38][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n47 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[38][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[39][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[39][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[40][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n49 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[40][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[41][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n50 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[41][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[42][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[42][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[43][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n52 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[43][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[44][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[44][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[45][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n54 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[45][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[46][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[46][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[47][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n56 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[47][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[48][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[48][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[49][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n58 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[49][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[50][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[50][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[51][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n60 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[51][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[52][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[52][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[53][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n62 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[53][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[54][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[54][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[55][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n64 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[55][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[56][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[56][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[57][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n66 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[57][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[58][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n67 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[58][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[59][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[59][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[60][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n69 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[60][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[61][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[61][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[62][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n71 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[62][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[63][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[63][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[24][3]  ( .D(\i_fifo_tx/n6 ), .E(\i_fifo_tx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[24][3] ) );
  DFEC1 \i_fifo_tx/mem_reg[0][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n10 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[0][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[1][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n11 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[1][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[2][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[2][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[3][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n13 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[3][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[4][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n14 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[4][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[5][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n15 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[5][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[6][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n16 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[6][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[7][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n17 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[7][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[8][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n18 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[8][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[9][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n19 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[9][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[10][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n20 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[10][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[11][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n21 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[11][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[12][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n22 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[12][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[13][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n23 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[13][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[14][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[14][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[15][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n25 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[15][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[16][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n26 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[16][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[17][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[17][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[18][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n28 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[18][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[19][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n29 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[19][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[20][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[20][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[21][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n31 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[21][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[22][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n32 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[22][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[23][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[23][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[25][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n34 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[25][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[26][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n35 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[26][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[27][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[27][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[28][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n37 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[28][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[29][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n38 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[29][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[30][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[30][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[31][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n40 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[31][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[32][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n41 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[32][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[33][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[33][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[34][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n43 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[34][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[35][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n44 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[35][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[36][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n45 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[36][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[37][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n46 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[37][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[38][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n47 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[38][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[39][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[39][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[40][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n49 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[40][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[41][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n50 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[41][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[42][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[42][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[43][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n52 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[43][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[44][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[44][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[45][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n54 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[45][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[46][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[46][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[47][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n56 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[47][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[48][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[48][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[49][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n58 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[49][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[50][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[50][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[51][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n60 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[51][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[52][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[52][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[53][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n62 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[53][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[54][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[54][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[55][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n64 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[55][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[56][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[56][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[57][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n66 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[57][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[58][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n67 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[58][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[59][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[59][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[60][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n69 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[60][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[61][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[61][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[62][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n71 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[62][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[63][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[63][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[24][4]  ( .D(\i_fifo_tx/n7 ), .E(\i_fifo_tx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[24][4] ) );
  DFEC1 \i_fifo_tx/mem_reg[0][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n10 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[0][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[1][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n11 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[1][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[2][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[2][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[3][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n13 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[3][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[4][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n14 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[4][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[5][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n15 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[5][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[6][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n16 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[6][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[7][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n17 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[7][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[8][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n18 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[8][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[9][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n19 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[9][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[10][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n20 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[10][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[11][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n21 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[11][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[12][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n22 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[12][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[13][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n23 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[13][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[14][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[14][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[15][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n25 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[15][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[16][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n26 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[16][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[17][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[17][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[18][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n28 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[18][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[19][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n29 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[19][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[20][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[20][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[21][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n31 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[21][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[22][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n32 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[22][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[23][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[23][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[25][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n34 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[25][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[26][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n35 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[26][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[27][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[27][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[28][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n37 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[28][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[29][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n38 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[29][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[30][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[30][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[31][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n40 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[31][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[32][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n41 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[32][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[33][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[33][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[34][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n43 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[34][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[35][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n44 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[35][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[36][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n45 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[36][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[37][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n46 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[37][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[38][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n47 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[38][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[39][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[39][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[40][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n49 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[40][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[41][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n50 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[41][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[42][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[42][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[43][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n52 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[43][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[44][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[44][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[45][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n54 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[45][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[46][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[46][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[47][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n56 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[47][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[48][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[48][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[49][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n58 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[49][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[50][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[50][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[51][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n60 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[51][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[52][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[52][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[53][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n62 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[53][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[54][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[54][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[55][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n64 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[55][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[56][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[56][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[57][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n66 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[57][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[58][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n67 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[58][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[59][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[59][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[60][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n69 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[60][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[61][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[61][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[62][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n71 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[62][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[63][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[63][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[24][5]  ( .D(\i_fifo_tx/n8 ), .E(\i_fifo_tx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[24][5] ) );
  DFEC1 \i_fifo_tx/mem_reg[0][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n10 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[0][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[1][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n11 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[1][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[2][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[2][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[3][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n13 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[3][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[4][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n14 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[4][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[5][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n15 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[5][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[6][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n16 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[6][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[7][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n17 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[7][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[8][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n18 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[8][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[9][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n19 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[9][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[10][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n20 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[10][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[11][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n21 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[11][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[12][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n22 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[12][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[13][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n23 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[13][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[14][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[14][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[15][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n25 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[15][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[16][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n26 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[16][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[17][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[17][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[18][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n28 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[18][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[19][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n29 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[19][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[20][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[20][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[21][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n31 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[21][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[22][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n32 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[22][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[23][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[23][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[25][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n34 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[25][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[26][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n35 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[26][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[27][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[27][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[28][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n37 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[28][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[29][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n38 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[29][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[30][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[30][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[31][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n40 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[31][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[32][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n41 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[32][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[33][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[33][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[34][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n43 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[34][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[35][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n44 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[35][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[36][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n45 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[36][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[37][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n46 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[37][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[38][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n47 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[38][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[39][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[39][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[40][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n49 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[40][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[41][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n50 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[41][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[42][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[42][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[43][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n52 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[43][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[44][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[44][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[45][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n54 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[45][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[46][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[46][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[47][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n56 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[47][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[48][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[48][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[49][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n58 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[49][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[50][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[50][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[51][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n60 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[51][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[52][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[52][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[53][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n62 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[53][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[54][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[54][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[55][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n64 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[55][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[56][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[56][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[57][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n66 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[57][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[58][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n67 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[58][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[59][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[59][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[60][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n69 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[60][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[61][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[61][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[62][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n71 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[62][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[63][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[63][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[24][6]  ( .D(\i_fifo_tx/n9 ), .E(\i_fifo_tx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[24][6] ) );
  DFEC1 \i_fifo_tx/mem_reg[0][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n10 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[0][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[1][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n11 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[1][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[2][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[2][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[3][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n13 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[3][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[4][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n14 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[4][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[5][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n15 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[5][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[6][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n16 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[6][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[7][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n17 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[7][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[8][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n18 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[8][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[9][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n19 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[9][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[10][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n20 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[10][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[11][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n21 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[11][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[12][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n22 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[12][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[13][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n23 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[13][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[14][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[14][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[15][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n25 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[15][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[16][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n26 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[16][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[17][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[17][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[18][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n28 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[18][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[19][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n29 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[19][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[20][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[20][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[21][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n31 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[21][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[22][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n32 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[22][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[23][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[23][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[25][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n34 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[25][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[26][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n35 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[26][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[27][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[27][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[28][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n37 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[28][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[29][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n38 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[29][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[30][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[30][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[31][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n40 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[31][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[32][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n41 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[32][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[33][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[33][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[34][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n43 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[34][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[35][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n44 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[35][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[36][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n45 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[36][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[37][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n46 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[37][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[38][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n47 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[38][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[39][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[39][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[40][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n49 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[40][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[41][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n50 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[41][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[42][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[42][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[43][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n52 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[43][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[44][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[44][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[45][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n54 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[45][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[46][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[46][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[47][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n56 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[47][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[48][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[48][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[49][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n58 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[49][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[50][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[50][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[51][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n60 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[51][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[52][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[52][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[53][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n62 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[53][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[54][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[54][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[55][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n64 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[55][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[56][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[56][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[57][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n66 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[57][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[58][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n67 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[58][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[59][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[59][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[60][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n69 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[60][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[61][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[61][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[62][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n71 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[62][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[63][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[63][7] ) );
  DFEC1 \i_fifo_tx/mem_reg[24][7]  ( .D(\i_fifo_tx/n73 ), .E(\i_fifo_tx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/mem[24][7] ) );
  DFEC1 \i_fifo_tx/rd_ptr_reg[1]  ( .D(\i_fifo_tx/N156 ), .E(\i_fifo_tx/n187 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/N31 ) );
  DFC1 \i_fifo_tx/compteur_reg[2]  ( .D(\i_fifo_tx/n206 ), .C(clk_i), .RN(
        resetn_i), .Q(\i_fifo_tx/N38 ) );
  DFC3 \i_fifo_tx/compteur_reg[1]  ( .D(\i_fifo_tx/n205 ), .C(clk_i), .RN(
        resetn_i), .Q(\i_fifo_tx/N37 ), .QN(\i_fifo_tx/n83 ) );
  DFC1 \i_fifo_tx/compteur_reg[0]  ( .D(\i_fifo_tx/n207 ), .C(clk_i), .RN(
        resetn_i), .Q(\i_fifo_tx/N36 ), .QN(\i_fifo_tx/n195 ) );
  CLKIN0 \i_cordic/U26  ( .A(\i_cordic/n22 ), .Q(\i_cordic/cor_x_s0[0][0] ) );
  AOI220 \i_cordic/U25  ( .A(\i_cordic/N14 ), .B(\i_cordic/S0/N32 ), .C(
        \i_cordic/ibb_ibuff [1]), .D(\i_cordic/n5 ), .Q(\i_cordic/n21 ) );
  AOI220 \i_cordic/U23  ( .A(\i_cordic/N15 ), .B(\i_cordic/S0/N32 ), .C(
        \i_cordic/ibb_ibuff [2]), .D(\i_cordic/n5 ), .Q(\i_cordic/n20 ) );
  AOI220 \i_cordic/U21  ( .A(\i_cordic/N16 ), .B(\i_cordic/S0/N32 ), .C(
        \i_cordic/ibb_ibuff [3]), .D(\i_cordic/n5 ), .Q(\i_cordic/n19 ) );
  NOR40 \i_cordic/U5  ( .A(\i_cordic/qbb_ibuff [3]), .B(
        \i_cordic/qbb_ibuff [2]), .C(\i_cordic/qbb_ibuff [1]), .D(
        \i_cordic/N6 ), .Q(\i_cordic/n6 ) );
  NAND20 \i_cordic/U4  ( .A(\i_cordic/qbb_ibuff [4]), .B(\i_cordic/n5 ), .Q(
        \i_cordic/n7 ) );
  DFC1 \i_cordic/wout_obuff_reg[5]  ( .D(\i_cordic/cor_w_s1[4][5] ), .C(clk_i), 
        .RN(resetn_i), .Q(cordic_phase_o[5]), .QN(n258) );
  DFC1 \i_cordic/wout_obuff_reg[4]  ( .D(\i_cordic/cor_w_s1[4][4] ), .C(clk_i), 
        .RN(resetn_i), .Q(cordic_phase_o[4]), .QN(n257) );
  DFC1 \i_cordic/wout_obuff_reg[3]  ( .D(\i_cordic/cor_w_s1[4][3] ), .C(clk_i), 
        .RN(resetn_i), .Q(cordic_phase_o[3]), .QN(n256) );
  DFC1 \i_cordic/wout_obuff_reg[2]  ( .D(\i_cordic/cor_w_s1[4][2] ), .C(clk_i), 
        .RN(resetn_i), .Q(cordic_phase_o[2]), .QN(n255) );
  DFC1 \i_cordic/wout_obuff_reg[1]  ( .D(\i_cordic/S2/n21 ), .C(clk_i), .RN(
        resetn_i), .Q(cordic_phase_o[1]), .QN(n254) );
  DFC1 \i_cordic/wout_obuff_reg[0]  ( .D(\*Logic1* ), .C(clk_i), .RN(resetn_i), 
        .Q(cordic_phase_o[0]), .QN(n253) );
  DFC1 \i_cordic/oValid_obuff_reg  ( .D(\i_cordic/valid_s1[4] ), .C(clk_i), 
        .RN(resetn_i), .Q(cordic_valid_o), .QN(n251) );
  DFC1 \i_cordic/cor_w_s1_reg[2][2]  ( .D(\*Logic1* ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/S2/N29 ), .QN(n117) );
  DFC1 \i_cordic/cor_w_s1_reg[2][3]  ( .D(\i_cordic/S1/sub_50/B_not [5]), .C(
        clk_i), .RN(resetn_i), .Q(\i_cordic/S2/N30 ) );
  DFC1 \i_cordic/cor_w_s1_reg[2][4]  ( .D(\i_cordic/cor_w_s0[2][4] ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/S2/N31 ), .QN(n101) );
  DFC1 \i_cordic/cor_w_s1_reg[2][5]  ( .D(\i_cordic/cor_w_s0[2][5] ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/S2/N32 ) );
  DFC1 \i_cordic/cor_y_s1_reg[2][0]  ( .D(\i_cordic/cor_y_s0[2][0] ), .C(clk_i), .RN(resetn_i), .QN(n225) );
  DFC1 \i_cordic/cor_y_s1_reg[2][1]  ( .D(\i_cordic/cor_y_s0[2][1] ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/cor_y_s1[2][1] ), .QN(n99) );
  DFC1 \i_cordic/cor_y_s1_reg[2][2]  ( .D(\i_cordic/cor_y_s0[2][2] ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/cor_y_s1[2][2] ), .QN(n229) );
  DFC1 \i_cordic/cor_y_s1_reg[2][3]  ( .D(\i_cordic/cor_y_s0[2][3] ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/cor_y_s1[2][3] ) );
  DFC1 \i_cordic/cor_y_s1_reg[2][4]  ( .D(\i_cordic/cor_y_s0[2][4] ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/cor_y_s1[2][4] ), .QN(n236) );
  DFC1 \i_cordic/cor_y_s1_reg[2][5]  ( .D(\i_cordic/cor_y_s0[2][5] ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/cor_y_s1[2][5] ), .QN(n185) );
  DFC1 \i_cordic/cor_x_s1_reg[2][2]  ( .D(\i_cordic/cor_x_s0[2][2] ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/cor_x_s1[2][2] ), .QN(n100) );
  DFC1 \i_cordic/cor_x_s1_reg[2][3]  ( .D(\i_cordic/cor_x_s0[2][3] ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/cor_x_s1[2][3] ), .QN(n218) );
  DFC1 \i_cordic/cor_x_s1_reg[2][4]  ( .D(\i_cordic/cor_x_s0[2][4] ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/cor_x_s1[2][4] ) );
  DFC1 \i_cordic/cor_x_s1_reg[2][5]  ( .D(\i_cordic/cor_x_s0[2][5] ), .C(clk_i), .RN(resetn_i), .Q(\i_cordic/cor_x_s1[2][5] ), .QN(n226) );
  DFC1 \i_cordic/valid_s1_reg[2]  ( .D(\i_cordic/valid_s0[2] ), .C(clk_i), 
        .RN(resetn_i), .Q(\i_cordic/valid_s1[4] ) );
  DFC1 \i_cordic/qbb_ibuff_reg[0]  ( .D(cordic_qbb_i[0]), .C(clk_i), .RN(
        resetn_i), .Q(\i_cordic/N6 ), .QN(\i_cordic/n16 ) );
  DFC1 \i_cordic/qbb_ibuff_reg[1]  ( .D(cordic_qbb_i[1]), .C(clk_i), .RN(
        resetn_i), .Q(\i_cordic/qbb_ibuff [1]), .QN(\i_cordic/n14 ) );
  DFC1 \i_cordic/qbb_ibuff_reg[2]  ( .D(cordic_qbb_i[2]), .C(clk_i), .RN(
        resetn_i), .Q(\i_cordic/qbb_ibuff [2]), .QN(\i_cordic/n12 ) );
  DFC1 \i_cordic/qbb_ibuff_reg[3]  ( .D(cordic_qbb_i[3]), .C(clk_i), .RN(
        resetn_i), .Q(\i_cordic/qbb_ibuff [3]), .QN(\i_cordic/n10 ) );
  DFC1 \i_cordic/qbb_ibuff_reg[4]  ( .D(cordic_qbb_i[4]), .C(clk_i), .RN(
        resetn_i), .Q(\i_cordic/qbb_ibuff [4]) );
  DFC1 \i_cordic/ibb_ibuff_reg[0]  ( .D(cordic_ibb_i[0]), .C(clk_i), .RN(
        resetn_i), .Q(\i_cordic/N13 ), .QN(n179) );
  DFC1 \i_cordic/ibb_ibuff_reg[1]  ( .D(cordic_ibb_i[1]), .C(clk_i), .RN(
        resetn_i), .Q(\i_cordic/ibb_ibuff [1]), .QN(n213) );
  DFC1 \i_cordic/ibb_ibuff_reg[2]  ( .D(cordic_ibb_i[2]), .C(clk_i), .RN(
        resetn_i), .Q(\i_cordic/ibb_ibuff [2]), .QN(n178) );
  DFC1 \i_cordic/ibb_ibuff_reg[3]  ( .D(cordic_ibb_i[3]), .C(clk_i), .RN(
        resetn_i), .Q(\i_cordic/ibb_ibuff [3]), .QN(n177) );
  DFC1 \i_cordic/iValid_ibuff_reg  ( .D(cordic_valid_i), .C(clk_i), .RN(
        resetn_i), .Q(\i_cordic/valid_s0[2] ) );
  NOR20 \i_fifo_rx/U221  ( .A(\i_fifo_rx/n188 ), .B(\i_fifo_rx/i [0]), .Q(
        \i_fifo_rx/N61 ) );
  CLKIN0 \i_fifo_rx/U220  ( .A(\i_fifo_rx/N54 ), .Q(\i_fifo_rx/n214 ) );
  NOR20 \i_fifo_rx/U219  ( .A(\i_fifo_rx/n188 ), .B(\i_fifo_rx/n214 ), .Q(
        \i_fifo_rx/N62 ) );
  CLKIN0 \i_fifo_rx/U218  ( .A(\i_fifo_rx/N55 ), .Q(\i_fifo_rx/n213 ) );
  NOR20 \i_fifo_rx/U217  ( .A(\i_fifo_rx/n188 ), .B(\i_fifo_rx/n213 ), .Q(
        \i_fifo_rx/N63 ) );
  CLKIN0 \i_fifo_rx/U216  ( .A(\i_fifo_rx/N56 ), .Q(\i_fifo_rx/n212 ) );
  NOR20 \i_fifo_rx/U215  ( .A(\i_fifo_rx/n188 ), .B(\i_fifo_rx/n212 ), .Q(
        \i_fifo_rx/N64 ) );
  CLKIN0 \i_fifo_rx/U214  ( .A(\i_fifo_rx/N57 ), .Q(\i_fifo_rx/n211 ) );
  NOR20 \i_fifo_rx/U213  ( .A(\i_fifo_rx/n188 ), .B(\i_fifo_rx/n211 ), .Q(
        \i_fifo_rx/N65 ) );
  CLKIN0 \i_fifo_rx/U212  ( .A(\i_fifo_rx/N58 ), .Q(\i_fifo_rx/n210 ) );
  NOR20 \i_fifo_rx/U211  ( .A(\i_fifo_rx/n188 ), .B(\i_fifo_rx/n210 ), .Q(
        \i_fifo_rx/N66 ) );
  CLKIN0 \i_fifo_rx/U210  ( .A(\i_fifo_rx/N59 ), .Q(\i_fifo_rx/n209 ) );
  NOR20 \i_fifo_rx/U209  ( .A(\i_fifo_rx/n188 ), .B(\i_fifo_rx/n209 ), .Q(
        \i_fifo_rx/N67 ) );
  NOR20 \i_fifo_rx/U207  ( .A(\i_fifo_rx/n188 ), .B(n238), .Q(\i_fifo_rx/N68 )
         );
  XNR20 \i_fifo_rx/U206  ( .A(\i_fifo_rx/wr_ptr[6] ), .B(\i_fifo_rx/rd_ptr[6] ), .Q(\i_fifo_rx/n174 ) );
  NAND20 \i_fifo_rx/U205  ( .A(\i_fifo_rx/N46 ), .B(\i_fifo_rx/n174 ), .Q(
        \i_fifo_rx/n11 ) );
  NOR20 \i_fifo_rx/U201  ( .A(\i_fifo_rx/n172 ), .B(n298), .Q(\i_fifo_rx/N680 ) );
  NOR20 \i_fifo_rx/U199  ( .A(\i_fifo_rx/n172 ), .B(n297), .Q(\i_fifo_rx/N681 ) );
  NOR20 \i_fifo_rx/U197  ( .A(\i_fifo_rx/n172 ), .B(n296), .Q(\i_fifo_rx/N682 ) );
  NOR20 \i_fifo_rx/U195  ( .A(\i_fifo_rx/n172 ), .B(n295), .Q(\i_fifo_rx/N683 ) );
  NOR20 \i_fifo_rx/U193  ( .A(\i_fifo_rx/n172 ), .B(n294), .Q(\i_fifo_rx/N684 ) );
  NOR20 \i_fifo_rx/U191  ( .A(\i_fifo_rx/n172 ), .B(n293), .Q(\i_fifo_rx/N685 ) );
  NOR20 \i_fifo_rx/U189  ( .A(\i_fifo_rx/n172 ), .B(n292), .Q(\i_fifo_rx/N686 ) );
  NOR20 \i_fifo_rx/U187  ( .A(\i_fifo_rx/n172 ), .B(n291), .Q(\i_fifo_rx/N687 ) );
  CLKIN0 \i_fifo_rx/U167  ( .A(\i_fifo_rx/N46 ), .Q(\i_fifo_rx/n175 ) );
  NAND20 \i_fifo_rx/U162  ( .A(\i_fifo_rx/n152 ), .B(\i_fifo_rx/n44 ), .Q(
        \i_fifo_rx/n169 ) );
  NAND20 \i_fifo_rx/U151  ( .A(\i_fifo_rx/n152 ), .B(\i_fifo_rx/n41 ), .Q(
        \i_fifo_rx/n167 ) );
  NAND20 \i_fifo_rx/U148  ( .A(\i_fifo_rx/n152 ), .B(\i_fifo_rx/n38 ), .Q(
        \i_fifo_rx/n165 ) );
  NAND20 \i_fifo_rx/U145  ( .A(\i_fifo_rx/n152 ), .B(\i_fifo_rx/n35 ), .Q(
        \i_fifo_rx/n163 ) );
  NAND20 \i_fifo_rx/U142  ( .A(\i_fifo_rx/n152 ), .B(\i_fifo_rx/n32 ), .Q(
        \i_fifo_rx/n161 ) );
  NAND20 \i_fifo_rx/U139  ( .A(\i_fifo_rx/n152 ), .B(\i_fifo_rx/n29 ), .Q(
        \i_fifo_rx/n159 ) );
  NAND20 \i_fifo_rx/U136  ( .A(\i_fifo_rx/n152 ), .B(\i_fifo_rx/n26 ), .Q(
        \i_fifo_rx/n157 ) );
  NAND20 \i_fifo_rx/U133  ( .A(\i_fifo_rx/n152 ), .B(\i_fifo_rx/n23 ), .Q(
        \i_fifo_rx/n151 ) );
  NAND20 \i_fifo_rx/U130  ( .A(\i_fifo_rx/n135 ), .B(\i_fifo_rx/n44 ), .Q(
        \i_fifo_rx/n149 ) );
  NAND20 \i_fifo_rx/U128  ( .A(\i_fifo_rx/n135 ), .B(\i_fifo_rx/n41 ), .Q(
        \i_fifo_rx/n147 ) );
  NAND20 \i_fifo_rx/U126  ( .A(\i_fifo_rx/n135 ), .B(\i_fifo_rx/n38 ), .Q(
        \i_fifo_rx/n145 ) );
  NAND20 \i_fifo_rx/U124  ( .A(\i_fifo_rx/n135 ), .B(\i_fifo_rx/n35 ), .Q(
        \i_fifo_rx/n143 ) );
  NAND20 \i_fifo_rx/U122  ( .A(\i_fifo_rx/n135 ), .B(\i_fifo_rx/n32 ), .Q(
        \i_fifo_rx/n141 ) );
  NAND20 \i_fifo_rx/U120  ( .A(\i_fifo_rx/n135 ), .B(\i_fifo_rx/n29 ), .Q(
        \i_fifo_rx/n139 ) );
  NAND20 \i_fifo_rx/U118  ( .A(\i_fifo_rx/n135 ), .B(\i_fifo_rx/n26 ), .Q(
        \i_fifo_rx/n137 ) );
  NAND20 \i_fifo_rx/U116  ( .A(\i_fifo_rx/n135 ), .B(\i_fifo_rx/n23 ), .Q(
        \i_fifo_rx/n134 ) );
  NAND20 \i_fifo_rx/U113  ( .A(\i_fifo_rx/n118 ), .B(\i_fifo_rx/n44 ), .Q(
        \i_fifo_rx/n132 ) );
  NAND20 \i_fifo_rx/U111  ( .A(\i_fifo_rx/n118 ), .B(\i_fifo_rx/n41 ), .Q(
        \i_fifo_rx/n130 ) );
  NAND20 \i_fifo_rx/U109  ( .A(\i_fifo_rx/n118 ), .B(\i_fifo_rx/n38 ), .Q(
        \i_fifo_rx/n128 ) );
  NAND20 \i_fifo_rx/U107  ( .A(\i_fifo_rx/n118 ), .B(\i_fifo_rx/n35 ), .Q(
        \i_fifo_rx/n126 ) );
  NAND20 \i_fifo_rx/U105  ( .A(\i_fifo_rx/n118 ), .B(\i_fifo_rx/n32 ), .Q(
        \i_fifo_rx/n124 ) );
  NAND20 \i_fifo_rx/U103  ( .A(\i_fifo_rx/n118 ), .B(\i_fifo_rx/n29 ), .Q(
        \i_fifo_rx/n122 ) );
  NAND20 \i_fifo_rx/U101  ( .A(\i_fifo_rx/n118 ), .B(\i_fifo_rx/n26 ), .Q(
        \i_fifo_rx/n120 ) );
  NAND20 \i_fifo_rx/U99  ( .A(\i_fifo_rx/n118 ), .B(\i_fifo_rx/n23 ), .Q(
        \i_fifo_rx/n117 ) );
  NAND20 \i_fifo_rx/U96  ( .A(\i_fifo_rx/n101 ), .B(\i_fifo_rx/n44 ), .Q(
        \i_fifo_rx/n115 ) );
  NAND20 \i_fifo_rx/U94  ( .A(\i_fifo_rx/n101 ), .B(\i_fifo_rx/n41 ), .Q(
        \i_fifo_rx/n113 ) );
  NAND20 \i_fifo_rx/U92  ( .A(\i_fifo_rx/n101 ), .B(\i_fifo_rx/n38 ), .Q(
        \i_fifo_rx/n111 ) );
  NAND20 \i_fifo_rx/U90  ( .A(\i_fifo_rx/n101 ), .B(\i_fifo_rx/n35 ), .Q(
        \i_fifo_rx/n109 ) );
  NAND20 \i_fifo_rx/U88  ( .A(\i_fifo_rx/n101 ), .B(\i_fifo_rx/n32 ), .Q(
        \i_fifo_rx/n107 ) );
  NAND20 \i_fifo_rx/U86  ( .A(\i_fifo_rx/n101 ), .B(\i_fifo_rx/n29 ), .Q(
        \i_fifo_rx/n105 ) );
  NAND20 \i_fifo_rx/U84  ( .A(\i_fifo_rx/n101 ), .B(\i_fifo_rx/n26 ), .Q(
        \i_fifo_rx/n103 ) );
  NAND20 \i_fifo_rx/U82  ( .A(\i_fifo_rx/n101 ), .B(\i_fifo_rx/n23 ), .Q(
        \i_fifo_rx/n100 ) );
  NAND20 \i_fifo_rx/U79  ( .A(\i_fifo_rx/n84 ), .B(\i_fifo_rx/n44 ), .Q(
        \i_fifo_rx/n98 ) );
  NAND20 \i_fifo_rx/U77  ( .A(\i_fifo_rx/n84 ), .B(\i_fifo_rx/n41 ), .Q(
        \i_fifo_rx/n96 ) );
  NAND20 \i_fifo_rx/U75  ( .A(\i_fifo_rx/n84 ), .B(\i_fifo_rx/n38 ), .Q(
        \i_fifo_rx/n94 ) );
  NAND20 \i_fifo_rx/U73  ( .A(\i_fifo_rx/n84 ), .B(\i_fifo_rx/n35 ), .Q(
        \i_fifo_rx/n92 ) );
  NAND20 \i_fifo_rx/U71  ( .A(\i_fifo_rx/n84 ), .B(\i_fifo_rx/n32 ), .Q(
        \i_fifo_rx/n90 ) );
  NAND20 \i_fifo_rx/U69  ( .A(\i_fifo_rx/n84 ), .B(\i_fifo_rx/n29 ), .Q(
        \i_fifo_rx/n88 ) );
  NAND20 \i_fifo_rx/U67  ( .A(\i_fifo_rx/n84 ), .B(\i_fifo_rx/n26 ), .Q(
        \i_fifo_rx/n86 ) );
  NAND20 \i_fifo_rx/U65  ( .A(\i_fifo_rx/n84 ), .B(\i_fifo_rx/n23 ), .Q(
        \i_fifo_rx/n83 ) );
  NAND20 \i_fifo_rx/U62  ( .A(\i_fifo_rx/n67 ), .B(\i_fifo_rx/n44 ), .Q(
        \i_fifo_rx/n81 ) );
  NAND20 \i_fifo_rx/U60  ( .A(\i_fifo_rx/n67 ), .B(\i_fifo_rx/n41 ), .Q(
        \i_fifo_rx/n79 ) );
  NAND20 \i_fifo_rx/U58  ( .A(\i_fifo_rx/n67 ), .B(\i_fifo_rx/n38 ), .Q(
        \i_fifo_rx/n77 ) );
  NAND20 \i_fifo_rx/U56  ( .A(\i_fifo_rx/n67 ), .B(\i_fifo_rx/n35 ), .Q(
        \i_fifo_rx/n75 ) );
  NAND20 \i_fifo_rx/U54  ( .A(\i_fifo_rx/n67 ), .B(\i_fifo_rx/n32 ), .Q(
        \i_fifo_rx/n73 ) );
  NAND20 \i_fifo_rx/U52  ( .A(\i_fifo_rx/n67 ), .B(\i_fifo_rx/n29 ), .Q(
        \i_fifo_rx/n71 ) );
  NAND20 \i_fifo_rx/U50  ( .A(\i_fifo_rx/n67 ), .B(\i_fifo_rx/n26 ), .Q(
        \i_fifo_rx/n69 ) );
  NAND20 \i_fifo_rx/U48  ( .A(\i_fifo_rx/n67 ), .B(\i_fifo_rx/n23 ), .Q(
        \i_fifo_rx/n66 ) );
  NAND20 \i_fifo_rx/U45  ( .A(\i_fifo_rx/n50 ), .B(\i_fifo_rx/n44 ), .Q(
        \i_fifo_rx/n64 ) );
  NAND20 \i_fifo_rx/U43  ( .A(\i_fifo_rx/n50 ), .B(\i_fifo_rx/n41 ), .Q(
        \i_fifo_rx/n62 ) );
  NAND20 \i_fifo_rx/U41  ( .A(\i_fifo_rx/n50 ), .B(\i_fifo_rx/n38 ), .Q(
        \i_fifo_rx/n60 ) );
  NAND20 \i_fifo_rx/U39  ( .A(\i_fifo_rx/n50 ), .B(\i_fifo_rx/n35 ), .Q(
        \i_fifo_rx/n58 ) );
  NAND20 \i_fifo_rx/U37  ( .A(\i_fifo_rx/n50 ), .B(\i_fifo_rx/n32 ), .Q(
        \i_fifo_rx/n56 ) );
  NAND20 \i_fifo_rx/U35  ( .A(\i_fifo_rx/n50 ), .B(\i_fifo_rx/n29 ), .Q(
        \i_fifo_rx/n54 ) );
  NAND20 \i_fifo_rx/U33  ( .A(\i_fifo_rx/n50 ), .B(\i_fifo_rx/n26 ), .Q(
        \i_fifo_rx/n52 ) );
  NAND20 \i_fifo_rx/U31  ( .A(\i_fifo_rx/n50 ), .B(\i_fifo_rx/n23 ), .Q(
        \i_fifo_rx/n49 ) );
  NAND20 \i_fifo_rx/U28  ( .A(\i_fifo_rx/n44 ), .B(\i_fifo_rx/n22 ), .Q(
        \i_fifo_rx/n43 ) );
  NAND20 \i_fifo_rx/U26  ( .A(\i_fifo_rx/n41 ), .B(\i_fifo_rx/n22 ), .Q(
        \i_fifo_rx/n40 ) );
  NAND20 \i_fifo_rx/U24  ( .A(\i_fifo_rx/n38 ), .B(\i_fifo_rx/n22 ), .Q(
        \i_fifo_rx/n37 ) );
  NAND20 \i_fifo_rx/U22  ( .A(\i_fifo_rx/n35 ), .B(\i_fifo_rx/n22 ), .Q(
        \i_fifo_rx/n34 ) );
  NAND20 \i_fifo_rx/U20  ( .A(\i_fifo_rx/n32 ), .B(\i_fifo_rx/n22 ), .Q(
        \i_fifo_rx/n31 ) );
  NAND20 \i_fifo_rx/U18  ( .A(\i_fifo_rx/n29 ), .B(\i_fifo_rx/n22 ), .Q(
        \i_fifo_rx/n28 ) );
  NAND20 \i_fifo_rx/U16  ( .A(\i_fifo_rx/n26 ), .B(\i_fifo_rx/n22 ), .Q(
        \i_fifo_rx/n25 ) );
  NAND20 \i_fifo_rx/U14  ( .A(\i_fifo_rx/n22 ), .B(\i_fifo_rx/n23 ), .Q(
        \i_fifo_rx/n14 ) );
  CLKIN0 \i_fifo_rx/U12  ( .A(\i_fifo_rx/n11 ), .Q(fifo_rx_pslv_err_o) );
  DF1 \i_fifo_rx/prdata_reg[0]  ( .D(\i_fifo_rx/N680 ), .C(clk_i), .Q(
        fifo_rx_prdata_o[0]) );
  DF1 \i_fifo_rx/prdata_reg[1]  ( .D(\i_fifo_rx/N681 ), .C(clk_i), .Q(
        fifo_rx_prdata_o[1]) );
  DF1 \i_fifo_rx/prdata_reg[2]  ( .D(\i_fifo_rx/N682 ), .C(clk_i), .Q(
        fifo_rx_prdata_o[2]) );
  DF1 \i_fifo_rx/prdata_reg[3]  ( .D(\i_fifo_rx/N683 ), .C(clk_i), .Q(
        fifo_rx_prdata_o[3]) );
  DF1 \i_fifo_rx/prdata_reg[4]  ( .D(\i_fifo_rx/N684 ), .C(clk_i), .Q(
        fifo_rx_prdata_o[4]) );
  DF1 \i_fifo_rx/prdata_reg[5]  ( .D(\i_fifo_rx/N685 ), .C(clk_i), .Q(
        fifo_rx_prdata_o[5]) );
  DF1 \i_fifo_rx/prdata_reg[6]  ( .D(\i_fifo_rx/N686 ), .C(clk_i), .Q(
        fifo_rx_prdata_o[6]) );
  DF1 \i_fifo_rx/prdata_reg[7]  ( .D(\i_fifo_rx/N687 ), .C(clk_i), .Q(
        fifo_rx_prdata_o[7]) );
  DFEC1 \i_fifo_rx/rd_ptr_reg[4]  ( .D(\i_fifo_rx/N692 ), .E(\i_fifo_rx/n173 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/N43 ) );
  DFEC1 \i_fifo_rx/rd_ptr_reg[6]  ( .D(\i_fifo_rx/N694 ), .E(\i_fifo_rx/n173 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/rd_ptr[6] ) );
  DFEC1 \i_fifo_rx/wr_ptr_reg[6]  ( .D(\i_fifo_rx/N86 ), .E(\i_fifo_rx/n171 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/wr_ptr[6] ) );
  DFE1 \i_fifo_rx/en_cdr_prec_reg  ( .D(fifo_rx_valid_i), .E(resetn_i), .C(
        clk_i), .QN(\i_fifo_rx/n176 ) );
  DFEC1 \i_fifo_rx/shift_register_reg[0]  ( .D(fifo_rx_data_i), .E(
        \i_fifo_rx/n177 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_fifo_rx/shift_register [0]) );
  DFEC1 \i_fifo_rx/shift_register_reg[1]  ( .D(fifo_rx_data_i), .E(
        \i_fifo_rx/n182 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_fifo_rx/shift_register [1]) );
  DFEC1 \i_fifo_rx/shift_register_reg[2]  ( .D(fifo_rx_data_i), .E(
        \i_fifo_rx/n184 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_fifo_rx/shift_register [2]) );
  DFEC1 \i_fifo_rx/shift_register_reg[3]  ( .D(fifo_rx_data_i), .E(
        \i_fifo_rx/n186 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_fifo_rx/shift_register [3]) );
  DFEC1 \i_fifo_rx/shift_register_reg[4]  ( .D(fifo_rx_data_i), .E(
        \i_fifo_rx/n189 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_fifo_rx/shift_register [4]) );
  DFEC1 \i_fifo_rx/shift_register_reg[5]  ( .D(fifo_rx_data_i), .E(
        \i_fifo_rx/n192 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_fifo_rx/shift_register [5]) );
  DFEC1 \i_fifo_rx/shift_register_reg[6]  ( .D(fifo_rx_data_i), .E(
        \i_fifo_rx/n194 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_fifo_rx/shift_register [6]) );
  DFEC1 \i_fifo_rx/shift_register_reg[7]  ( .D(fifo_rx_data_i), .E(
        \i_fifo_rx/n196 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_fifo_rx/shift_register [7]) );
  DFC1 \i_fifo_rx/i_reg[1]  ( .D(\i_fifo_rx/N62 ), .C(clk_i), .RN(resetn_i), 
        .Q(\i_fifo_rx/i [1]), .QN(\i_fifo_rx/n180 ) );
  DFC1 \i_fifo_rx/i_reg[2]  ( .D(\i_fifo_rx/N63 ), .C(clk_i), .RN(resetn_i), 
        .Q(\i_fifo_rx/i [2]), .QN(\i_fifo_rx/n198 ) );
  DFC1 \i_fifo_rx/i_reg[3]  ( .D(\i_fifo_rx/N64 ), .C(clk_i), .RN(resetn_i), 
        .Q(\i_fifo_rx/i [3]), .QN(n105) );
  DFC1 \i_fifo_rx/i_reg[4]  ( .D(\i_fifo_rx/N65 ), .C(clk_i), .RN(resetn_i), 
        .Q(\i_fifo_rx/i [4]), .QN(n104) );
  DFC1 \i_fifo_rx/i_reg[5]  ( .D(\i_fifo_rx/N66 ), .C(clk_i), .RN(resetn_i), 
        .Q(\i_fifo_rx/i [5]) );
  DFC1 \i_fifo_rx/i_reg[6]  ( .D(\i_fifo_rx/N67 ), .C(clk_i), .RN(resetn_i), 
        .Q(\i_fifo_rx/i [6]) );
  DFC1 \i_fifo_rx/i_reg[7]  ( .D(\i_fifo_rx/N68 ), .C(clk_i), .RN(resetn_i), 
        .Q(\i_fifo_rx/i [7]) );
  DFC1 \i_fifo_rx/i_reg[0]  ( .D(\i_fifo_rx/N61 ), .C(clk_i), .RN(resetn_i), 
        .Q(\i_fifo_rx/i [0]), .QN(\i_fifo_rx/n179 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U192  ( .A(mod_iq_enable_i), .Q(
        \i_mod_iq/fsm_mapping/n214 ) );
  NOR20 \i_mod_iq/fsm_mapping/U191  ( .A(\i_mod_iq/fsm_mapping/n214 ), .B(
        \i_mod_iq/fsm_mapping/en_prev ), .Q(\i_mod_iq/fsm_mapping/N260 ) );
  NOR20 \i_mod_iq/fsm_mapping/U190  ( .A(\i_mod_iq/fsm_mapping/C_STATE [1]), 
        .B(\i_mod_iq/fsm_mapping/C_STATE [0]), .Q(\i_mod_iq/fsm_mapping/n127 )
         );
  CLKIN0 \i_mod_iq/fsm_mapping/U189  ( .A(\i_mod_iq/fsm_mapping/n127 ), .Q(
        \i_mod_iq/fsm_mapping/n116 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U187  ( .A(fifo_tx_mem_state_o), .Q(
        \i_mod_iq/fsm_mapping/n215 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U185  ( .A(\i_mod_iq/fsm_mapping/n173 ), .Q(
        \i_mod_iq/fsm_mapping/n115 ) );
  NOR30 \i_mod_iq/fsm_mapping/U184  ( .A(\i_mod_iq/fsm_mapping/cpt [0]), .B(
        \i_mod_iq/fsm_mapping/cpt [1]), .C(\i_mod_iq/fsm_mapping/n69 ), .Q(
        \i_mod_iq/fsm_mapping/n217 ) );
  NOR30 \i_mod_iq/fsm_mapping/U183  ( .A(\i_mod_iq/fsm_mapping/cpt_old [0]), 
        .B(\i_mod_iq/fsm_mapping/cpt_old [1]), .C(\i_mod_iq/fsm_mapping/n218 ), 
        .Q(\i_mod_iq/fsm_mapping/n216 ) );
  NAND30 \i_mod_iq/fsm_mapping/U182  ( .A(\i_mod_iq/fsm_mapping/n217 ), .B(
        \i_mod_iq/fsm_mapping/n215 ), .C(\i_mod_iq/fsm_mapping/n216 ), .Q(
        \i_mod_iq/fsm_mapping/n208 ) );
  NAND20 \i_mod_iq/fsm_mapping/U178  ( .A(\i_mod_iq/fsm_mapping/n51 ), .B(
        \i_mod_iq/fsm_mapping/n90 ), .Q(\i_mod_iq/fsm_mapping/n188 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U177  ( .A(\i_mod_iq/fsm_mapping/n217 ), .Q(
        \i_mod_iq/fsm_mapping/n180 ) );
  NOR20 \i_mod_iq/fsm_mapping/U176  ( .A(\i_mod_iq/fsm_mapping/n214 ), .B(
        \i_mod_iq/fsm_mapping/n180 ), .Q(\i_mod_iq/fsm_mapping/n120 ) );
  NAND20 \i_mod_iq/fsm_mapping/U175  ( .A(\i_mod_iq/fsm_mapping/n216 ), .B(
        \i_mod_iq/fsm_mapping/n120 ), .Q(\i_mod_iq/fsm_mapping/n210 ) );
  NAND20 \i_mod_iq/fsm_mapping/U172  ( .A(\i_mod_iq/fsm_mapping/n69 ), .B(
        \i_mod_iq/fsm_mapping/n98 ), .Q(\i_mod_iq/fsm_mapping/n83 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U171  ( .A(\i_mod_iq/fsm_mapping/n83 ), .Q(
        \i_mod_iq/fsm_mapping/n195 ) );
  NOR30 \i_mod_iq/fsm_mapping/U169  ( .A(\i_mod_iq/fsm_mapping/cpt_old [1]), 
        .B(\i_mod_iq/fsm_mapping/cpt_old [2]), .C(\i_mod_iq/fsm_mapping/n80 ), 
        .Q(\i_mod_iq/fsm_mapping/n161 ) );
  NAND30 \i_mod_iq/fsm_mapping/U168  ( .A(\i_mod_iq/fsm_mapping/n179 ), .B(
        \i_mod_iq/fsm_mapping/n215 ), .C(\i_mod_iq/fsm_mapping/n161 ), .Q(
        \i_mod_iq/fsm_mapping/n207 ) );
  NOR20 \i_mod_iq/fsm_mapping/U167  ( .A(\i_mod_iq/fsm_mapping/n80 ), .B(
        \i_mod_iq/fsm_mapping/n214 ), .Q(\i_mod_iq/fsm_mapping/n143 ) );
  NAND30 \i_mod_iq/fsm_mapping/U166  ( .A(\i_mod_iq/fsm_mapping/n119 ), .B(
        \i_mod_iq/fsm_mapping/n207 ), .C(\i_mod_iq/fsm_mapping/n143 ), .Q(
        \i_mod_iq/fsm_mapping/n213 ) );
  NOR40 \i_mod_iq/fsm_mapping/U165  ( .A(\i_mod_iq/fsm_mapping/n213 ), .B(
        \i_mod_iq/fsm_mapping/cpt_old [0]), .C(
        \i_mod_iq/fsm_mapping/cpt_old [2]), .D(
        \i_mod_iq/fsm_mapping/cpt_old [1]), .Q(\i_mod_iq/fsm_mapping/n212 ) );
  AOI310 \i_mod_iq/fsm_mapping/U164  ( .A(\i_mod_iq/fsm_mapping/n208 ), .B(
        \i_mod_iq/fsm_mapping/n188 ), .C(\i_mod_iq/fsm_mapping/n210 ), .D(
        \i_mod_iq/fsm_mapping/n212 ), .Q(\i_mod_iq/fsm_mapping/n211 ) );
  OAI310 \i_mod_iq/fsm_mapping/U163  ( .A(\i_mod_iq/fsm_mapping/n116 ), .B(
        \i_mod_iq/fsm_mapping/en_prev ), .C(\i_mod_iq/fsm_mapping/n115 ), .D(
        \i_mod_iq/fsm_mapping/n211 ), .Q(\i_mod_iq/fsm_mapping/N_STATE [0]) );
  OAI210 \i_mod_iq/fsm_mapping/U162  ( .A(\i_mod_iq/fsm_mapping/n210 ), .B(
        \i_mod_iq/fsm_mapping/n51 ), .C(\i_mod_iq/fsm_mapping/n90 ), .Q(
        \i_mod_iq/fsm_mapping/n209 ) );
  AOI220 \i_mod_iq/fsm_mapping/U161  ( .A(\i_mod_iq/fsm_mapping/n207 ), .B(
        \i_mod_iq/fsm_mapping/n119 ), .C(\i_mod_iq/fsm_mapping/n208 ), .D(
        \i_mod_iq/fsm_mapping/n209 ), .Q(\i_mod_iq/fsm_mapping/n206 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U160  ( .A(\i_mod_iq/fsm_mapping/n206 ), .Q(
        \i_mod_iq/fsm_mapping/N_STATE [1]) );
  NOR20 \i_mod_iq/fsm_mapping/U159  ( .A(\i_mod_iq/fsm_mapping/n98 ), .B(
        \i_mod_iq/fsm_mapping/n163 ), .Q(\i_mod_iq/fsm_mapping/n205 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U158  ( .A(\i_mod_iq/fsm_mapping/n188 ), .Q(
        \i_mod_iq/fsm_mapping/n204 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U156  ( .A(\i_mod_iq/fsm_mapping/n90 ), .Q(
        \i_mod_iq/fsm_mapping/n47 ) );
  OAI210 \i_mod_iq/fsm_mapping/U154  ( .A(\i_mod_iq/fsm_mapping/n205 ), .B(
        \i_mod_iq/fsm_mapping/n204 ), .C(\i_mod_iq/fsm_mapping/n193 ), .Q(
        \i_mod_iq/fsm_mapping/n201 ) );
  NAND20 \i_mod_iq/fsm_mapping/U153  ( .A(\i_mod_iq/fsm_mapping/n205 ), .B(
        \i_mod_iq/fsm_mapping/n69 ), .Q(\i_mod_iq/fsm_mapping/n154 ) );
  NOR20 \i_mod_iq/fsm_mapping/U152  ( .A(\i_mod_iq/fsm_mapping/n204 ), .B(
        \i_mod_iq/fsm_mapping/n154 ), .Q(\i_mod_iq/fsm_mapping/n202 ) );
  XNR20 \i_mod_iq/fsm_mapping/U151  ( .A(\i_mod_iq/fsm_mapping/cpt [1]), .B(
        \i_mod_iq/fsm_mapping/cpt [0]), .Q(\i_mod_iq/fsm_mapping/n82 ) );
  AOI2110 \i_mod_iq/fsm_mapping/U150  ( .A(\i_mod_iq/fsm_mapping/n82 ), .B(
        \i_mod_iq/fsm_mapping/n98 ), .C(\i_mod_iq/fsm_mapping/n53 ), .D(
        \i_mod_iq/fsm_mapping/n69 ), .Q(\i_mod_iq/fsm_mapping/n203 ) );
  AOI2110 \i_mod_iq/fsm_mapping/U149  ( .A(\i_mod_iq/fsm_mapping/cpt [2]), .B(
        \i_mod_iq/fsm_mapping/n201 ), .C(\i_mod_iq/fsm_mapping/n202 ), .D(
        \i_mod_iq/fsm_mapping/n203 ), .Q(\i_mod_iq/fsm_mapping/n196 ) );
  NOR20 \i_mod_iq/fsm_mapping/U147  ( .A(n252), .B(\i_mod_iq/fsm_mapping/n164 ), .Q(\i_mod_iq/fsm_mapping/n197 ) );
  NOR20 \i_mod_iq/fsm_mapping/U146  ( .A(\i_mod_iq/fsm_mapping/n68 ), .B(
        \i_mod_iq/fsm_mapping/n119 ), .Q(\i_mod_iq/fsm_mapping/n174 ) );
  OAI210 \i_mod_iq/fsm_mapping/U145  ( .A(\i_mod_iq/fsm_mapping/C_STATE [0]), 
        .B(\i_mod_iq/fsm_mapping/n173 ), .C(\i_mod_iq/fsm_mapping/n174 ), .Q(
        \i_mod_iq/fsm_mapping/n199 ) );
  OAI210 \i_mod_iq/fsm_mapping/U140  ( .A(\i_mod_iq/fsm_mapping/n197 ), .B(
        \i_mod_iq/fsm_mapping/n199 ), .C(\i_mod_iq/fsm_mapping/N259 ), .Q(
        \i_mod_iq/fsm_mapping/n182 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U139  ( .A(\i_mod_iq/fsm_mapping/n182 ), .Q(
        \i_mod_iq/fsm_mapping/n183 ) );
  NAND20 \i_mod_iq/fsm_mapping/U138  ( .A(\i_mod_iq/fsm_mapping/n119 ), .B(
        \i_mod_iq/fsm_mapping/n80 ), .Q(\i_mod_iq/fsm_mapping/n65 ) );
  AOI220 \i_mod_iq/fsm_mapping/U136  ( .A(\i_mod_iq/fsm_mapping/n194 ), .B(
        \i_mod_iq/fsm_mapping/n98 ), .C(\i_mod_iq/fsm_mapping/n195 ), .D(
        \i_mod_iq/fsm_mapping/n188 ), .Q(\i_mod_iq/fsm_mapping/n191 ) );
  NOR20 \i_mod_iq/fsm_mapping/U135  ( .A(\i_mod_iq/fsm_mapping/n69 ), .B(
        \i_mod_iq/fsm_mapping/n193 ), .Q(\i_mod_iq/fsm_mapping/n184 ) );
  OAI210 \i_mod_iq/fsm_mapping/U134  ( .A(\i_mod_iq/fsm_mapping/n184 ), .B(
        \i_mod_iq/fsm_mapping/n182 ), .C(\i_mod_iq/fsm_mapping/cpt [0]), .Q(
        \i_mod_iq/fsm_mapping/n192 ) );
  OAI210 \i_mod_iq/fsm_mapping/U133  ( .A(\i_mod_iq/fsm_mapping/n191 ), .B(
        \i_mod_iq/fsm_mapping/n182 ), .C(\i_mod_iq/fsm_mapping/n192 ), .Q(
        \i_mod_iq/fsm_mapping/n232 ) );
  AOI210 \i_mod_iq/fsm_mapping/U128  ( .A(\i_mod_iq/fsm_mapping/n184 ), .B(
        \i_mod_iq/fsm_mapping/cpt [1]), .C(\i_mod_iq/fsm_mapping/n185 ), .Q(
        \i_mod_iq/fsm_mapping/n181 ) );
  NOR40 \i_mod_iq/fsm_mapping/U127  ( .A(\i_mod_iq/fsm_mapping/n178 ), .B(
        \i_mod_iq/fsm_mapping/n179 ), .C(\i_mod_iq/fsm_mapping/n180 ), .D(
        \i_mod_iq/fsm_mapping/cpt_old [2]), .Q(\i_mod_iq/fsm_mapping/n166 ) );
  XNR20 \i_mod_iq/fsm_mapping/U125  ( .A(\i_mod_iq/fsm_mapping/b_in_prev ), 
        .B(mod_iq_data_i), .Q(\i_mod_iq/fsm_mapping/n114 ) );
  NAND20 \i_mod_iq/fsm_mapping/U124  ( .A(\i_mod_iq/fsm_mapping/n143 ), .B(
        \i_mod_iq/fsm_mapping/n114 ), .Q(\i_mod_iq/fsm_mapping/n170 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U123  ( .A(\i_mod_iq/fsm_mapping/n170 ), .Q(
        \i_mod_iq/fsm_mapping/n175 ) );
  OAI210 \i_mod_iq/fsm_mapping/U121  ( .A(\i_mod_iq/fsm_mapping/C_STATE [1]), 
        .B(\i_mod_iq/fsm_mapping/n173 ), .C(\i_mod_iq/fsm_mapping/n174 ), .Q(
        \i_mod_iq/fsm_mapping/n171 ) );
  NOR20 \i_mod_iq/fsm_mapping/U119  ( .A(\i_mod_iq/fsm_mapping/n170 ), .B(
        \i_mod_iq/fsm_mapping/n168 ), .Q(\i_mod_iq/fsm_mapping/n169 ) );
  OAI220 \i_mod_iq/fsm_mapping/U118  ( .A(\i_mod_iq/fsm_mapping/n167 ), .B(
        \i_mod_iq/fsm_mapping/n168 ), .C(\i_mod_iq/fsm_mapping/n169 ), .D(
        \i_mod_iq/fsm_mapping/n131 ), .Q(\i_mod_iq/fsm_mapping/n230 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U117  ( .A(\i_mod_iq/fsm_mapping/n120 ), .Q(
        \i_mod_iq/fsm_mapping/n113 ) );
  NAND20 \i_mod_iq/fsm_mapping/U116  ( .A(\i_mod_iq/fsm_mapping/n166 ), .B(
        \i_mod_iq/fsm_mapping/n113 ), .Q(\i_mod_iq/fsm_mapping/n75 ) );
  NAND20 \i_mod_iq/fsm_mapping/U115  ( .A(\i_mod_iq/fsm_mapping/cpt [2]), .B(
        \i_mod_iq/fsm_mapping/n75 ), .Q(\i_mod_iq/fsm_mapping/n58 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U114  ( .A(\i_mod_iq/fsm_mapping/n58 ), .Q(
        \i_mod_iq/fsm_mapping/n59 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U112  ( .A(\i_mod_iq/fsm_mapping/n44 ), .Q(
        \i_mod_iq/fsm_mapping/n45 ) );
  NAND20 \i_mod_iq/fsm_mapping/U111  ( .A(\i_mod_iq/fsm_mapping/n69 ), .B(
        \i_mod_iq/fsm_mapping/n163 ), .Q(\i_mod_iq/fsm_mapping/n99 ) );
  OAI2110 \i_mod_iq/fsm_mapping/U108  ( .A(\i_mod_iq/fsm_mapping/n69 ), .B(
        \i_mod_iq/fsm_mapping/n156 ), .C(\i_mod_iq/fsm_mapping/n75 ), .D(
        \i_mod_iq/fsm_mapping/n81 ), .Q(\i_mod_iq/fsm_mapping/n157 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U107  ( .A(\i_mod_iq/fsm_mapping/n80 ), .Q(
        \i_mod_iq/fsm_mapping/n56 ) );
  NAND20 \i_mod_iq/fsm_mapping/U106  ( .A(\i_mod_iq/fsm_mapping/n161 ), .B(
        \i_mod_iq/fsm_mapping/cpt_old [0]), .Q(\i_mod_iq/fsm_mapping/n145 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U101  ( .A(\i_mod_iq/fsm_mapping/n92 ), .Q(
        \i_mod_iq/fsm_mapping/n54 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U99  ( .A(\i_mod_iq/fsm_mapping/n154 ), .Q(
        \i_mod_iq/fsm_mapping/n160 ) );
  OAI220 \i_mod_iq/fsm_mapping/U98  ( .A(\i_mod_iq/fsm_mapping/n159 ), .B(
        \i_mod_iq/fsm_mapping/n53 ), .C(\i_mod_iq/fsm_mapping/n160 ), .D(
        \i_mod_iq/fsm_mapping/n90 ), .Q(\i_mod_iq/fsm_mapping/n158 ) );
  AOI210 \i_mod_iq/fsm_mapping/U97  ( .A(\i_mod_iq/fsm_mapping/n68 ), .B(
        \i_mod_iq/fsm_mapping/n157 ), .C(\i_mod_iq/fsm_mapping/n158 ), .Q(
        \i_mod_iq/fsm_mapping/n155 ) );
  NAND20 \i_mod_iq/fsm_mapping/U96  ( .A(\i_mod_iq/fsm_mapping/n154 ), .B(
        \i_mod_iq/fsm_mapping/n83 ), .Q(\i_mod_iq/fsm_mapping/n153 ) );
  AOI220 \i_mod_iq/fsm_mapping/U95  ( .A(\i_mod_iq/fsm_mapping/n153 ), .B(
        \i_mod_iq/fsm_mapping/n131 ), .C(\i_mod_iq/fsm_mapping/S_AQ ), .D(
        \i_mod_iq/fsm_mapping/n83 ), .Q(\i_mod_iq/fsm_mapping/n151 ) );
  NOR20 \i_mod_iq/fsm_mapping/U93  ( .A(\i_mod_iq/fsm_mapping/n69 ), .B(
        \i_mod_iq/fsm_mapping/n147 ), .Q(\i_mod_iq/fsm_mapping/n152 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U92  ( .A(\i_mod_iq/fsm_mapping/n75 ), .Q(
        \i_mod_iq/fsm_mapping/n138 ) );
  AOI2110 \i_mod_iq/fsm_mapping/U91  ( .A(\i_mod_iq/fsm_mapping/cpt [0]), .B(
        \i_mod_iq/fsm_mapping/n69 ), .C(\i_mod_iq/fsm_mapping/n152 ), .D(
        \i_mod_iq/fsm_mapping/n138 ), .Q(\i_mod_iq/fsm_mapping/n150 ) );
  OAI220 \i_mod_iq/fsm_mapping/U90  ( .A(\i_mod_iq/fsm_mapping/n150 ), .B(
        \i_mod_iq/fsm_mapping/n51 ), .C(\i_mod_iq/fsm_mapping/n151 ), .D(
        \i_mod_iq/fsm_mapping/n90 ), .Q(\i_mod_iq/fsm_mapping/n149 ) );
  AOI210 \i_mod_iq/fsm_mapping/U89  ( .A(\i_mod_iq/fsm_mapping/n119 ), .B(
        \i_mod_iq/fsm_mapping/n148 ), .C(\i_mod_iq/fsm_mapping/n149 ), .Q(
        \i_mod_iq/fsm_mapping/n146 ) );
  XNR20 \i_mod_iq/fsm_mapping/U88  ( .A(\i_mod_iq/fsm_mapping/n131 ), .B(
        \i_mod_iq/fsm_mapping/n99 ), .Q(\i_mod_iq/fsm_mapping/n139 ) );
  OAI220 \i_mod_iq/fsm_mapping/U83  ( .A(\i_mod_iq/fsm_mapping/n76 ), .B(
        \i_mod_iq/fsm_mapping/n134 ), .C(\i_mod_iq/fsm_mapping/n139 ), .D(
        \i_mod_iq/fsm_mapping/n90 ), .Q(\i_mod_iq/fsm_mapping/n136 ) );
  AOI210 \i_mod_iq/fsm_mapping/U82  ( .A(\i_mod_iq/fsm_mapping/n69 ), .B(
        \i_mod_iq/fsm_mapping/cpt [1]), .C(\i_mod_iq/fsm_mapping/n138 ), .Q(
        \i_mod_iq/fsm_mapping/n106 ) );
  AOI2110 \i_mod_iq/fsm_mapping/U80  ( .A(\i_mod_iq/fsm_mapping/n119 ), .B(
        \i_mod_iq/fsm_mapping/n135 ), .C(\i_mod_iq/fsm_mapping/n136 ), .D(
        \i_mod_iq/fsm_mapping/n137 ), .Q(\i_mod_iq/fsm_mapping/n133 ) );
  AOI210 \i_mod_iq/fsm_mapping/U79  ( .A(\i_mod_iq/fsm_mapping/n68 ), .B(
        \i_mod_iq/fsm_mapping/n59 ), .C(\i_mod_iq/fsm_mapping/n45 ), .Q(
        \i_mod_iq/fsm_mapping/n128 ) );
  AOI220 \i_mod_iq/fsm_mapping/U77  ( .A(\i_mod_iq/fsm_mapping/n47 ), .B(
        \i_mod_iq/fsm_mapping/n131 ), .C(\i_mod_iq/fsm_mapping/n119 ), .D(
        \i_mod_iq/fsm_mapping/n132 ), .Q(\i_mod_iq/fsm_mapping/n130 ) );
  OAI220 \i_mod_iq/fsm_mapping/U76  ( .A(\i_mod_iq/fsm_mapping/n128 ), .B(
        \i_mod_iq/fsm_mapping/n129 ), .C(\i_mod_iq/fsm_mapping/n45 ), .D(
        \i_mod_iq/fsm_mapping/n130 ), .Q(\i_mod_iq/fsm_mapping/n229 ) );
  AOI220 \i_mod_iq/fsm_mapping/U73  ( .A(\i_mod_iq/fsm_mapping/temp_QBB [0]), 
        .B(\i_mod_iq/fsm_mapping/n39 ), .C(mod_iq_qbb_o[0]), .D(
        \i_mod_iq/fsm_mapping/n40 ), .Q(\i_mod_iq/fsm_mapping/n126 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U72  ( .A(\i_mod_iq/fsm_mapping/n126 ), .Q(
        \i_mod_iq/fsm_mapping/n228 ) );
  AOI220 \i_mod_iq/fsm_mapping/U71  ( .A(\i_mod_iq/fsm_mapping/temp_QBB [1]), 
        .B(\i_mod_iq/fsm_mapping/n39 ), .C(mod_iq_qbb_o[1]), .D(
        \i_mod_iq/fsm_mapping/n40 ), .Q(\i_mod_iq/fsm_mapping/n125 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U70  ( .A(\i_mod_iq/fsm_mapping/n125 ), .Q(
        \i_mod_iq/fsm_mapping/n227 ) );
  AOI220 \i_mod_iq/fsm_mapping/U69  ( .A(\i_mod_iq/fsm_mapping/temp_QBB [2]), 
        .B(\i_mod_iq/fsm_mapping/n39 ), .C(mod_iq_qbb_o[2]), .D(
        \i_mod_iq/fsm_mapping/n40 ), .Q(\i_mod_iq/fsm_mapping/n124 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U68  ( .A(\i_mod_iq/fsm_mapping/n124 ), .Q(
        \i_mod_iq/fsm_mapping/n226 ) );
  AOI220 \i_mod_iq/fsm_mapping/U67  ( .A(\i_mod_iq/fsm_mapping/temp_QBB [3]), 
        .B(\i_mod_iq/fsm_mapping/n39 ), .C(mod_iq_qbb_o[3]), .D(
        \i_mod_iq/fsm_mapping/n40 ), .Q(\i_mod_iq/fsm_mapping/n123 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U66  ( .A(\i_mod_iq/fsm_mapping/n123 ), .Q(
        \i_mod_iq/fsm_mapping/n225 ) );
  NAND20 \i_mod_iq/fsm_mapping/U64  ( .A(\i_mod_iq/fsm_mapping/n120 ), .B(n192), .Q(\i_mod_iq/fsm_mapping/n118 ) );
  AOI210 \i_mod_iq/fsm_mapping/U63  ( .A(\i_mod_iq/fsm_mapping/n47 ), .B(
        \i_mod_iq/fsm_mapping/n118 ), .C(\i_mod_iq/fsm_mapping/n119 ), .Q(
        \i_mod_iq/fsm_mapping/n117 ) );
  AOI210 \i_mod_iq/fsm_mapping/U61  ( .A(\i_mod_iq/fsm_mapping/n68 ), .B(
        \i_mod_iq/fsm_mapping/n113 ), .C(\i_mod_iq/fsm_mapping/n109 ), .Q(
        \i_mod_iq/fsm_mapping/n107 ) );
  NOR20 \i_mod_iq/fsm_mapping/U60  ( .A(\i_mod_iq/fsm_mapping/n115 ), .B(
        \i_mod_iq/fsm_mapping/n116 ), .Q(\i_mod_iq/fsm_mapping/n110 ) );
  XNR20 \i_mod_iq/fsm_mapping/U59  ( .A(\i_mod_iq/fsm_mapping/n48 ), .B(
        \i_mod_iq/fsm_mapping/n114 ), .Q(\i_mod_iq/fsm_mapping/n111 ) );
  OAI210 \i_mod_iq/fsm_mapping/U58  ( .A(\i_mod_iq/fsm_mapping/n76 ), .B(
        \i_mod_iq/fsm_mapping/n113 ), .C(\i_mod_iq/fsm_mapping/n90 ), .Q(
        \i_mod_iq/fsm_mapping/n112 ) );
  AOI220 \i_mod_iq/fsm_mapping/U57  ( .A(\i_mod_iq/fsm_mapping/n110 ), .B(
        mod_iq_data_i), .C(\i_mod_iq/fsm_mapping/n111 ), .D(
        \i_mod_iq/fsm_mapping/n112 ), .Q(\i_mod_iq/fsm_mapping/n108 ) );
  OAI220 \i_mod_iq/fsm_mapping/U56  ( .A(\i_mod_iq/fsm_mapping/n107 ), .B(
        \i_mod_iq/fsm_mapping/n48 ), .C(\i_mod_iq/fsm_mapping/n108 ), .D(
        \i_mod_iq/fsm_mapping/n109 ), .Q(\i_mod_iq/fsm_mapping/n224 ) );
  OAI2110 \i_mod_iq/fsm_mapping/U55  ( .A(\i_mod_iq/fsm_mapping/n100 ), .B(
        \i_mod_iq/fsm_mapping/n58 ), .C(\i_mod_iq/fsm_mapping/n83 ), .D(
        \i_mod_iq/fsm_mapping/n106 ), .Q(\i_mod_iq/fsm_mapping/n102 ) );
  NOR20 \i_mod_iq/fsm_mapping/U54  ( .A(\i_mod_iq/fsm_mapping/n99 ), .B(
        \i_mod_iq/fsm_mapping/n98 ), .Q(\i_mod_iq/fsm_mapping/n105 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U53  ( .A(\i_mod_iq/fsm_mapping/n105 ), .Q(
        \i_mod_iq/fsm_mapping/n97 ) );
  AOI220 \i_mod_iq/fsm_mapping/U52  ( .A(\i_mod_iq/fsm_mapping/n54 ), .B(
        \i_mod_iq/fsm_mapping/temp_IBB [0]), .C(\i_mod_iq/fsm_mapping/n92 ), 
        .D(\i_mod_iq/fsm_mapping/n97 ), .Q(\i_mod_iq/fsm_mapping/n104 ) );
  OAI220 \i_mod_iq/fsm_mapping/U51  ( .A(\i_mod_iq/fsm_mapping/n104 ), .B(
        \i_mod_iq/fsm_mapping/n53 ), .C(\i_mod_iq/fsm_mapping/n105 ), .D(
        \i_mod_iq/fsm_mapping/n90 ), .Q(\i_mod_iq/fsm_mapping/n103 ) );
  AOI210 \i_mod_iq/fsm_mapping/U50  ( .A(\i_mod_iq/fsm_mapping/n68 ), .B(
        \i_mod_iq/fsm_mapping/n102 ), .C(\i_mod_iq/fsm_mapping/n103 ), .Q(
        \i_mod_iq/fsm_mapping/n101 ) );
  OAI210 \i_mod_iq/fsm_mapping/U49  ( .A(\i_mod_iq/fsm_mapping/n59 ), .B(
        \i_mod_iq/fsm_mapping/n98 ), .C(\i_mod_iq/fsm_mapping/n99 ), .Q(
        \i_mod_iq/fsm_mapping/n96 ) );
  NAND20 \i_mod_iq/fsm_mapping/U48  ( .A(\i_mod_iq/fsm_mapping/n98 ), .B(
        \i_mod_iq/fsm_mapping/n99 ), .Q(\i_mod_iq/fsm_mapping/n93 ) );
  AOI210 \i_mod_iq/fsm_mapping/U47  ( .A(\i_mod_iq/fsm_mapping/n93 ), .B(
        \i_mod_iq/fsm_mapping/n97 ), .C(\i_mod_iq/fsm_mapping/S_AI ), .Q(
        \i_mod_iq/fsm_mapping/n94 ) );
  AOI220 \i_mod_iq/fsm_mapping/U46  ( .A(\i_mod_iq/fsm_mapping/S_AI ), .B(
        \i_mod_iq/fsm_mapping/n96 ), .C(\i_mod_iq/fsm_mapping/n94 ), .D(
        \i_mod_iq/fsm_mapping/n58 ), .Q(\i_mod_iq/fsm_mapping/n95 ) );
  OAI210 \i_mod_iq/fsm_mapping/U45  ( .A(\i_mod_iq/fsm_mapping/n84 ), .B(
        \i_mod_iq/fsm_mapping/n58 ), .C(\i_mod_iq/fsm_mapping/n95 ), .Q(
        \i_mod_iq/fsm_mapping/n86 ) );
  AOI210 \i_mod_iq/fsm_mapping/U44  ( .A(\i_mod_iq/fsm_mapping/S_AI ), .B(
        \i_mod_iq/fsm_mapping/n93 ), .C(\i_mod_iq/fsm_mapping/n94 ), .Q(
        \i_mod_iq/fsm_mapping/n89 ) );
  OAI220 \i_mod_iq/fsm_mapping/U41  ( .A(\i_mod_iq/fsm_mapping/n88 ), .B(
        \i_mod_iq/fsm_mapping/n53 ), .C(\i_mod_iq/fsm_mapping/n89 ), .D(
        \i_mod_iq/fsm_mapping/n90 ), .Q(\i_mod_iq/fsm_mapping/n87 ) );
  AOI210 \i_mod_iq/fsm_mapping/U40  ( .A(\i_mod_iq/fsm_mapping/n68 ), .B(
        \i_mod_iq/fsm_mapping/n86 ), .C(\i_mod_iq/fsm_mapping/n87 ), .Q(
        \i_mod_iq/fsm_mapping/n85 ) );
  NAND20 \i_mod_iq/fsm_mapping/U39  ( .A(\i_mod_iq/fsm_mapping/n82 ), .B(
        \i_mod_iq/fsm_mapping/n83 ), .Q(\i_mod_iq/fsm_mapping/n67 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U38  ( .A(\i_mod_iq/fsm_mapping/n67 ), .Q(
        \i_mod_iq/fsm_mapping/n77 ) );
  OAI220 \i_mod_iq/fsm_mapping/U37  ( .A(\i_mod_iq/fsm_mapping/n81 ), .B(
        \i_mod_iq/fsm_mapping/n51 ), .C(\i_mod_iq/fsm_mapping/n77 ), .D(
        \i_mod_iq/fsm_mapping/n65 ), .Q(\i_mod_iq/fsm_mapping/n62 ) );
  NOR20 \i_mod_iq/fsm_mapping/U35  ( .A(\i_mod_iq/fsm_mapping/n53 ), .B(
        \i_mod_iq/fsm_mapping/n80 ), .Q(\i_mod_iq/fsm_mapping/n73 ) );
  NOR20 \i_mod_iq/fsm_mapping/U34  ( .A(\i_mod_iq/fsm_mapping/n76 ), .B(
        \i_mod_iq/fsm_mapping/n75 ), .Q(\i_mod_iq/fsm_mapping/n79 ) );
  AOI2110 \i_mod_iq/fsm_mapping/U33  ( .A(n85), .B(\i_mod_iq/fsm_mapping/n73 ), 
        .C(\i_mod_iq/fsm_mapping/n79 ), .D(\i_mod_iq/fsm_mapping/n47 ), .Q(
        \i_mod_iq/fsm_mapping/n70 ) );
  XNR20 \i_mod_iq/fsm_mapping/U32  ( .A(\i_mod_iq/fsm_mapping/S_AI ), .B(
        \i_mod_iq/fsm_mapping/n77 ), .Q(\i_mod_iq/fsm_mapping/n71 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U31  ( .A(\i_mod_iq/fsm_mapping/n76 ), .Q(
        \i_mod_iq/fsm_mapping/n74 ) );
  AOI220 \i_mod_iq/fsm_mapping/U30  ( .A(\i_mod_iq/fsm_mapping/n73 ), .B(
        \i_mod_iq/fsm_mapping/n57 ), .C(\i_mod_iq/fsm_mapping/n74 ), .D(
        \i_mod_iq/fsm_mapping/n75 ), .Q(\i_mod_iq/fsm_mapping/n72 ) );
  OAI220 \i_mod_iq/fsm_mapping/U29  ( .A(\i_mod_iq/fsm_mapping/n70 ), .B(
        \i_mod_iq/fsm_mapping/n71 ), .C(\i_mod_iq/fsm_mapping/n72 ), .D(
        \i_mod_iq/fsm_mapping/n60 ), .Q(\i_mod_iq/fsm_mapping/n63 ) );
  NAND20 \i_mod_iq/fsm_mapping/U28  ( .A(\i_mod_iq/fsm_mapping/n68 ), .B(
        \i_mod_iq/fsm_mapping/n69 ), .Q(\i_mod_iq/fsm_mapping/n66 ) );
  AOI2110 \i_mod_iq/fsm_mapping/U27  ( .A(\i_mod_iq/fsm_mapping/n65 ), .B(
        \i_mod_iq/fsm_mapping/n66 ), .C(\i_mod_iq/fsm_mapping/n67 ), .D(
        \i_mod_iq/fsm_mapping/S_AI ), .Q(\i_mod_iq/fsm_mapping/n64 ) );
  AOI2110 \i_mod_iq/fsm_mapping/U26  ( .A(\i_mod_iq/fsm_mapping/S_AI ), .B(
        \i_mod_iq/fsm_mapping/n62 ), .C(\i_mod_iq/fsm_mapping/n63 ), .D(
        \i_mod_iq/fsm_mapping/n64 ), .Q(\i_mod_iq/fsm_mapping/n61 ) );
  AOI210 \i_mod_iq/fsm_mapping/U24  ( .A(\i_mod_iq/fsm_mapping/n56 ), .B(
        \i_mod_iq/fsm_mapping/n57 ), .C(\i_mod_iq/fsm_mapping/S_AI ), .Q(
        \i_mod_iq/fsm_mapping/n55 ) );
  AOI210 \i_mod_iq/fsm_mapping/U23  ( .A(\i_mod_iq/fsm_mapping/n54 ), .B(
        \i_mod_iq/fsm_mapping/temp_IBB [3]), .C(\i_mod_iq/fsm_mapping/n55 ), 
        .Q(\i_mod_iq/fsm_mapping/n52 ) );
  OAI220 \i_mod_iq/fsm_mapping/U22  ( .A(\i_mod_iq/fsm_mapping/n50 ), .B(
        \i_mod_iq/fsm_mapping/n51 ), .C(\i_mod_iq/fsm_mapping/n52 ), .D(
        \i_mod_iq/fsm_mapping/n53 ), .Q(\i_mod_iq/fsm_mapping/n49 ) );
  AOI210 \i_mod_iq/fsm_mapping/U21  ( .A(\i_mod_iq/fsm_mapping/n47 ), .B(
        \i_mod_iq/fsm_mapping/n48 ), .C(\i_mod_iq/fsm_mapping/n49 ), .Q(
        \i_mod_iq/fsm_mapping/n46 ) );
  AOI220 \i_mod_iq/fsm_mapping/U20  ( .A(\i_mod_iq/fsm_mapping/temp_IBB [0]), 
        .B(\i_mod_iq/fsm_mapping/n39 ), .C(mod_iq_ibb_o[0]), .D(
        \i_mod_iq/fsm_mapping/n40 ), .Q(\i_mod_iq/fsm_mapping/n43 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U19  ( .A(\i_mod_iq/fsm_mapping/n43 ), .Q(
        \i_mod_iq/fsm_mapping/n223 ) );
  AOI220 \i_mod_iq/fsm_mapping/U18  ( .A(\i_mod_iq/fsm_mapping/temp_IBB [1]), 
        .B(\i_mod_iq/fsm_mapping/n39 ), .C(mod_iq_ibb_o[1]), .D(
        \i_mod_iq/fsm_mapping/n40 ), .Q(\i_mod_iq/fsm_mapping/n42 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U17  ( .A(\i_mod_iq/fsm_mapping/n42 ), .Q(
        \i_mod_iq/fsm_mapping/n222 ) );
  AOI220 \i_mod_iq/fsm_mapping/U16  ( .A(\i_mod_iq/fsm_mapping/temp_IBB [2]), 
        .B(\i_mod_iq/fsm_mapping/n39 ), .C(mod_iq_ibb_o[2]), .D(
        \i_mod_iq/fsm_mapping/n40 ), .Q(\i_mod_iq/fsm_mapping/n41 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U15  ( .A(\i_mod_iq/fsm_mapping/n41 ), .Q(
        \i_mod_iq/fsm_mapping/n221 ) );
  AOI220 \i_mod_iq/fsm_mapping/U14  ( .A(\i_mod_iq/fsm_mapping/temp_IBB [3]), 
        .B(\i_mod_iq/fsm_mapping/n39 ), .C(mod_iq_ibb_o[3]), .D(
        \i_mod_iq/fsm_mapping/n40 ), .Q(\i_mod_iq/fsm_mapping/n38 ) );
  CLKIN0 \i_mod_iq/fsm_mapping/U13  ( .A(\i_mod_iq/fsm_mapping/n38 ), .Q(
        \i_mod_iq/fsm_mapping/n220 ) );
  INV2 \i_mod_iq/fsm_mapping/U12  ( .A(\i_mod_iq/fsm_mapping/n196 ), .Q(
        \i_mod_iq/fsm_mapping/n37 ) );
  INV2 \i_mod_iq/fsm_mapping/U11  ( .A(\i_mod_iq/fsm_mapping/N261 ), .Q(
        \i_mod_iq/fsm_mapping/n36 ) );
  INV2 \i_mod_iq/fsm_mapping/U10  ( .A(\i_mod_iq/fsm_mapping/n181 ), .Q(
        \i_mod_iq/fsm_mapping/n35 ) );
  INV2 \i_mod_iq/fsm_mapping/U9  ( .A(\i_mod_iq/fsm_mapping/n101 ), .Q(
        \i_mod_iq/fsm_mapping/n34 ) );
  INV2 \i_mod_iq/fsm_mapping/U8  ( .A(\i_mod_iq/fsm_mapping/n146 ), .Q(
        \i_mod_iq/fsm_mapping/n33 ) );
  INV2 \i_mod_iq/fsm_mapping/U7  ( .A(\i_mod_iq/fsm_mapping/n155 ), .Q(
        \i_mod_iq/fsm_mapping/n32 ) );
  INV2 \i_mod_iq/fsm_mapping/U6  ( .A(\i_mod_iq/fsm_mapping/n85 ), .Q(
        \i_mod_iq/fsm_mapping/n31 ) );
  INV2 \i_mod_iq/fsm_mapping/U5  ( .A(\i_mod_iq/fsm_mapping/n61 ), .Q(
        \i_mod_iq/fsm_mapping/n30 ) );
  INV2 \i_mod_iq/fsm_mapping/U4  ( .A(\i_mod_iq/fsm_mapping/n46 ), .Q(
        \i_mod_iq/fsm_mapping/n29 ) );
  INV2 \i_mod_iq/fsm_mapping/U3  ( .A(\i_mod_iq/fsm_mapping/n133 ), .Q(
        \i_mod_iq/fsm_mapping/n28 ) );
  DFC1 \i_mod_iq/fsm_mapping/QBB_reg[2]  ( .D(\i_mod_iq/fsm_mapping/n226 ), 
        .C(clk_i), .RN(resetn_i), .Q(mod_iq_qbb_o[2]) );
  DFEC1 \i_mod_iq/fsm_mapping/temp_QBB_reg[2]  ( .D(\i_mod_iq/fsm_mapping/n28 ), .E(\i_mod_iq/fsm_mapping/n44 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/temp_QBB [2]), .QN(\i_mod_iq/fsm_mapping/n134 )
         );
  DFC1 \i_mod_iq/fsm_mapping/IBB_reg[3]  ( .D(\i_mod_iq/fsm_mapping/n220 ), 
        .C(clk_i), .RN(resetn_i), .Q(mod_iq_ibb_o[3]) );
  DFEC1 \i_mod_iq/fsm_mapping/temp_IBB_reg[3]  ( .D(\i_mod_iq/fsm_mapping/n29 ), .E(\i_mod_iq/fsm_mapping/n44 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/temp_IBB [3]) );
  DFC1 \i_mod_iq/fsm_mapping/IBB_reg[2]  ( .D(\i_mod_iq/fsm_mapping/n221 ), 
        .C(clk_i), .RN(resetn_i), .Q(mod_iq_ibb_o[2]) );
  DFEC1 \i_mod_iq/fsm_mapping/temp_IBB_reg[2]  ( .D(\i_mod_iq/fsm_mapping/n30 ), .E(\i_mod_iq/fsm_mapping/n44 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/temp_IBB [2]), .QN(\i_mod_iq/fsm_mapping/n60 )
         );
  DFC1 \i_mod_iq/fsm_mapping/IBB_reg[1]  ( .D(\i_mod_iq/fsm_mapping/n222 ), 
        .C(clk_i), .RN(resetn_i), .Q(mod_iq_ibb_o[1]) );
  DFEC1 \i_mod_iq/fsm_mapping/temp_IBB_reg[1]  ( .D(\i_mod_iq/fsm_mapping/n31 ), .E(\i_mod_iq/fsm_mapping/n44 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/temp_IBB [1]), .QN(\i_mod_iq/fsm_mapping/n84 )
         );
  DFC1 \i_mod_iq/fsm_mapping/S_AI_reg  ( .D(\i_mod_iq/fsm_mapping/n224 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_mod_iq/fsm_mapping/S_AI ), .QN(
        \i_mod_iq/fsm_mapping/n48 ) );
  DFC1 \i_mod_iq/fsm_mapping/QBB_reg[0]  ( .D(\i_mod_iq/fsm_mapping/n228 ), 
        .C(clk_i), .RN(resetn_i), .Q(mod_iq_qbb_o[0]) );
  DFEC1 \i_mod_iq/fsm_mapping/temp_QBB_reg[0]  ( .D(\i_mod_iq/fsm_mapping/n32 ), .E(\i_mod_iq/fsm_mapping/n44 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/temp_QBB [0]), .QN(\i_mod_iq/fsm_mapping/n156 )
         );
  DFC1 \i_mod_iq/fsm_mapping/QBB_reg[1]  ( .D(\i_mod_iq/fsm_mapping/n227 ), 
        .C(clk_i), .RN(resetn_i), .Q(mod_iq_qbb_o[1]) );
  DFEC1 \i_mod_iq/fsm_mapping/temp_QBB_reg[1]  ( .D(\i_mod_iq/fsm_mapping/n33 ), .E(\i_mod_iq/fsm_mapping/n44 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/temp_QBB [1]), .QN(\i_mod_iq/fsm_mapping/n147 )
         );
  DFC1 \i_mod_iq/fsm_mapping/QBB_reg[3]  ( .D(\i_mod_iq/fsm_mapping/n225 ), 
        .C(clk_i), .RN(resetn_i), .Q(mod_iq_qbb_o[3]) );
  DFC1 \i_mod_iq/fsm_mapping/temp_QBB_reg[3]  ( .D(\i_mod_iq/fsm_mapping/n229 ), .C(clk_i), .RN(resetn_i), .Q(\i_mod_iq/fsm_mapping/temp_QBB [3]), .QN(
        \i_mod_iq/fsm_mapping/n129 ) );
  DFC1 \i_mod_iq/fsm_mapping/IBB_reg[0]  ( .D(\i_mod_iq/fsm_mapping/n223 ), 
        .C(clk_i), .RN(resetn_i), .Q(mod_iq_ibb_o[0]) );
  DFEC1 \i_mod_iq/fsm_mapping/temp_IBB_reg[0]  ( .D(\i_mod_iq/fsm_mapping/n34 ), .E(\i_mod_iq/fsm_mapping/n44 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/temp_IBB [0]), .QN(\i_mod_iq/fsm_mapping/n100 )
         );
  DFP1 \i_mod_iq/fsm_mapping/S_AQ_reg  ( .D(\i_mod_iq/fsm_mapping/n230 ), .C(
        clk_i), .SN(resetn_i), .Q(\i_mod_iq/fsm_mapping/S_AQ ), .QN(
        \i_mod_iq/fsm_mapping/n131 ) );
  DFEC1 \i_mod_iq/fsm_mapping/ready_reg  ( .D(\i_mod_iq/fsm_mapping/n177 ), 
        .E(\i_mod_iq/fsm_mapping/N259 ), .C(clk_i), .RN(resetn_i), .QN(n115)
         );
  DFP1 \i_mod_iq/fsm_mapping/f_dac_down_reg  ( .D(\i_mod_iq/fsm_mapping/n231 ), 
        .C(clk_i), .SN(resetn_i), .QN(\i_mod_iq/fsm_mapping/n177 ) );
  DFEC1 \i_mod_iq/fsm_mapping/cpt_reg[1]  ( .D(\i_mod_iq/fsm_mapping/n35 ), 
        .E(\i_mod_iq/fsm_mapping/n183 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/cpt [1]), .QN(\i_mod_iq/fsm_mapping/n163 ) );
  DFEC1 \i_mod_iq/fsm_mapping/cpt_old_reg[0]  ( .D(
        \i_mod_iq/fsm_mapping/cpt [0]), .E(\i_mod_iq/fsm_mapping/N259 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_mod_iq/fsm_mapping/cpt_old [0]), .QN(
        \i_mod_iq/fsm_mapping/n179 ) );
  DFC1 \i_mod_iq/fsm_mapping/cpt_reg[0]  ( .D(\i_mod_iq/fsm_mapping/n232 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_mod_iq/fsm_mapping/cpt [0]), .QN(
        \i_mod_iq/fsm_mapping/n98 ) );
  DFC1 \i_mod_iq/fsm_mapping/en_dac_reg  ( .D(\i_mod_iq/en_10MHz ), .C(clk_i), 
        .RN(\i_mod_iq/fsm_mapping/n36 ), .Q(mod_iq_valid_o) );
  DFC1 \i_mod_iq/fsm_mapping/C_STATE_reg[1]  ( .D(
        \i_mod_iq/fsm_mapping/N_STATE [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/C_STATE [1]) );
  DFEC1 \i_mod_iq/fsm_mapping/cpt_old_reg[2]  ( .D(
        \i_mod_iq/fsm_mapping/cpt [2]), .E(\i_mod_iq/fsm_mapping/N259 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_mod_iq/fsm_mapping/cpt_old [2]), .QN(
        \i_mod_iq/fsm_mapping/n218 ) );
  DFC1 \i_mod_iq/fsm_mapping/C_STATE_reg[0]  ( .D(
        \i_mod_iq/fsm_mapping/N_STATE [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/C_STATE [0]), .QN(\i_mod_iq/fsm_mapping/n164 )
         );
  DFEC1 \i_mod_iq/fsm_mapping/b_in_prev_reg  ( .D(
        \i_mod_iq/fsm_mapping/s_b_in_prev ), .E(\i_mod_iq/fsm_mapping/N259 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_mod_iq/fsm_mapping/b_in_prev ) );
  DFEC1 \i_mod_iq/fsm_mapping/s_b_in_prev_reg  ( .D(mod_iq_data_i), .E(
        \i_mod_iq/fsm_mapping/N260 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/s_b_in_prev ) );
  DFC1 \i_mod_iq/fsm_mapping/en_prev_reg  ( .D(mod_iq_enable_i), .C(clk_i), 
        .RN(resetn_i), .Q(\i_mod_iq/fsm_mapping/en_prev ) );
  DFC1 \i_mod_iq/fsm_mapping/en_10MHz_prev_reg  ( .D(\i_mod_iq/en_10MHz ), .C(
        clk_i), .RN(resetn_i), .Q(\i_mod_iq/fsm_mapping/en_10MHz_prev ) );
  DFC1 \i_mod_iq/fsm_mapping/dac_ready_prev_reg  ( .D(\*Logic1* ), .C(clk_i), 
        .RN(resetn_i), .Q(n192), .QN(n252) );
  NOR30 \i_mod_iq/en_gen_map/U7  ( .A(\i_mod_iq/en_gen_map/cpt [0]), .B(
        \i_mod_iq/en_gen_map/cpt [1]), .C(\i_mod_iq/en_gen_map/n3 ), .Q(
        \i_mod_iq/en_gen_map/N13 ) );
  NOR20 \i_mod_iq/en_gen_map/U6  ( .A(\i_mod_iq/en_gen_map/cpt [0]), .B(
        \i_mod_iq/en_gen_map/N13 ), .Q(\i_mod_iq/en_gen_map/N6 ) );
  XNR20 \i_mod_iq/en_gen_map/U5  ( .A(\i_mod_iq/en_gen_map/cpt [1]), .B(
        \i_mod_iq/en_gen_map/cpt [0]), .Q(\i_mod_iq/en_gen_map/n4 ) );
  DFC1 \i_mod_iq/en_gen_map/clk_out_reg  ( .D(\i_mod_iq/en_gen_map/N13 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_mod_iq/en_10MHz ), .QN(n237) );
  JKC1 \i_mod_iq/en_gen_map/cpt_reg[2]  ( .J(\i_mod_iq/en_gen_map/n1 ), .K(
        \i_mod_iq/en_gen_map/n4 ), .C(clk_i), .RN(resetn_i), .QN(
        \i_mod_iq/en_gen_map/n3 ) );
  TFEC1 \i_mod_iq/en_gen_map/cpt_reg[1]  ( .T(\i_mod_iq/en_gen_map/cpt [0]), 
        .C(clk_i), .RN(resetn_i), .Q(\i_mod_iq/en_gen_map/cpt [1]), .QN(n122)
         );
  DFC1 \i_mod_iq/en_gen_map/cpt_reg[0]  ( .D(\i_mod_iq/en_gen_map/N6 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_mod_iq/en_gen_map/cpt [0]), .QN(n123) );
  CLKIN0 \i_iq_demod/demod/U54  ( .A(\i_iq_demod/demod/N36 ), .Q(
        \i_iq_demod/demod/n43 ) );
  CLKIN0 \i_iq_demod/demod/U51  ( .A(demod_iq_iif_i[1]), .Q(
        \i_iq_demod/demod/n41 ) );
  OAI220 \i_iq_demod/demod/U50  ( .A(\i_iq_demod/demod/n32 ), .B(n282), .C(
        \i_iq_demod/demod/n33 ), .D(\i_iq_demod/demod/n41 ), .Q(
        \i_iq_demod/demod/IC [1]) );
  CLKIN0 \i_iq_demod/demod/U48  ( .A(demod_iq_iif_i[2]), .Q(
        \i_iq_demod/demod/n39 ) );
  OAI220 \i_iq_demod/demod/U47  ( .A(\i_iq_demod/demod/n32 ), .B(n283), .C(
        \i_iq_demod/demod/n33 ), .D(\i_iq_demod/demod/n39 ), .Q(
        \i_iq_demod/demod/IC [2]) );
  CLKIN0 \i_iq_demod/demod/U45  ( .A(demod_iq_iif_i[3]), .Q(
        \i_iq_demod/demod/n37 ) );
  OAI220 \i_iq_demod/demod/U44  ( .A(\i_iq_demod/demod/n32 ), .B(n284), .C(
        \i_iq_demod/demod/n33 ), .D(\i_iq_demod/demod/n37 ), .Q(
        \i_iq_demod/demod/IC [3]) );
  CLKIN0 \i_iq_demod/demod/U42  ( .A(demod_iq_iif_i[4]), .Q(
        \i_iq_demod/demod/n35 ) );
  OAI220 \i_iq_demod/demod/U41  ( .A(\i_iq_demod/demod/n32 ), .B(n285), .C(
        \i_iq_demod/demod/n33 ), .D(\i_iq_demod/demod/n35 ), .Q(
        \i_iq_demod/demod/IC [4]) );
  OAI220 \i_iq_demod/demod/U36  ( .A(\i_iq_demod/demod/n20 ), .B(n282), .C(
        \i_iq_demod/demod/n22 ), .D(\i_iq_demod/demod/n41 ), .Q(
        \i_iq_demod/demod/IS [1]) );
  OAI220 \i_iq_demod/demod/U35  ( .A(\i_iq_demod/demod/n20 ), .B(n283), .C(
        \i_iq_demod/demod/n22 ), .D(\i_iq_demod/demod/n39 ), .Q(
        \i_iq_demod/demod/IS [2]) );
  OAI220 \i_iq_demod/demod/U34  ( .A(\i_iq_demod/demod/n20 ), .B(n284), .C(
        \i_iq_demod/demod/n22 ), .D(\i_iq_demod/demod/n37 ), .Q(
        \i_iq_demod/demod/IS [3]) );
  OAI220 \i_iq_demod/demod/U33  ( .A(\i_iq_demod/demod/n20 ), .B(n285), .C(
        \i_iq_demod/demod/n22 ), .D(\i_iq_demod/demod/n35 ), .Q(
        \i_iq_demod/demod/IS [4]) );
  CLKIN0 \i_iq_demod/demod/U31  ( .A(\i_iq_demod/demod/N41 ), .Q(
        \i_iq_demod/demod/n31 ) );
  CLKIN0 \i_iq_demod/demod/U28  ( .A(demod_iq_qif_i[1]), .Q(
        \i_iq_demod/demod/n29 ) );
  OAI220 \i_iq_demod/demod/U27  ( .A(n281), .B(\i_iq_demod/demod/n32 ), .C(
        \i_iq_demod/demod/n29 ), .D(\i_iq_demod/demod/n33 ), .Q(
        \i_iq_demod/demod/QC [1]) );
  CLKIN0 \i_iq_demod/demod/U25  ( .A(demod_iq_qif_i[2]), .Q(
        \i_iq_demod/demod/n27 ) );
  OAI220 \i_iq_demod/demod/U24  ( .A(n280), .B(\i_iq_demod/demod/n32 ), .C(
        \i_iq_demod/demod/n27 ), .D(\i_iq_demod/demod/n33 ), .Q(
        \i_iq_demod/demod/QC [2]) );
  CLKIN0 \i_iq_demod/demod/U22  ( .A(demod_iq_qif_i[3]), .Q(
        \i_iq_demod/demod/n25 ) );
  OAI220 \i_iq_demod/demod/U21  ( .A(n279), .B(\i_iq_demod/demod/n32 ), .C(
        \i_iq_demod/demod/n25 ), .D(\i_iq_demod/demod/n33 ), .Q(
        \i_iq_demod/demod/QC [3]) );
  CLKIN0 \i_iq_demod/demod/U19  ( .A(demod_iq_qif_i[4]), .Q(
        \i_iq_demod/demod/n23 ) );
  OAI220 \i_iq_demod/demod/U18  ( .A(n278), .B(\i_iq_demod/demod/n32 ), .C(
        \i_iq_demod/demod/n23 ), .D(\i_iq_demod/demod/n33 ), .Q(
        \i_iq_demod/demod/QC [4]) );
  OAI220 \i_iq_demod/demod/U16  ( .A(\i_iq_demod/demod/n20 ), .B(n281), .C(
        \i_iq_demod/demod/n22 ), .D(\i_iq_demod/demod/n29 ), .Q(
        \i_iq_demod/demod/QS [1]) );
  OAI220 \i_iq_demod/demod/U15  ( .A(\i_iq_demod/demod/n20 ), .B(n280), .C(
        \i_iq_demod/demod/n22 ), .D(\i_iq_demod/demod/n27 ), .Q(
        \i_iq_demod/demod/QS [2]) );
  OAI220 \i_iq_demod/demod/U14  ( .A(\i_iq_demod/demod/n20 ), .B(n279), .C(
        \i_iq_demod/demod/n22 ), .D(\i_iq_demod/demod/n25 ), .Q(
        \i_iq_demod/demod/QS [3]) );
  OAI220 \i_iq_demod/demod/U13  ( .A(\i_iq_demod/demod/n20 ), .B(n278), .C(
        \i_iq_demod/demod/n22 ), .D(\i_iq_demod/demod/n23 ), .Q(
        \i_iq_demod/demod/QS [4]) );
  NOR20 \i_iq_demod/filtre_I/U95  ( .A(\i_iq_demod/filtre_I/shift_count [2]), 
        .B(\i_iq_demod/filtre_I/shift_count [0]), .Q(\i_iq_demod/filtre_I/n42 ) );
  NAND20 \i_iq_demod/filtre_I/U40  ( .A(\i_iq_demod/filtre_I/current_state [1]), .B(\i_iq_demod/filtre_I/n2 ), .Q(\i_iq_demod/filtre_I/n10 ) );
  OAI220 \i_iq_demod/filtre_I/U39  ( .A(\i_iq_demod/filtre_I/current_state [1]), .B(\i_iq_demod/filtre_I/next_state [0]), .C(\i_iq_demod/filtre_I/n10 ), .D(
        \i_iq_demod/filtre_I/current_state [0]), .Q(
        \i_iq_demod/filtre_I/next_state [1]) );
  CLKIN0 \i_iq_demod/filtre_I/U37  ( .A(\i_iq_demod/filtre_I/n10 ), .Q(
        \i_iq_demod/filtre_I/n7 ) );
  AOI210 \i_iq_demod/filtre_I/U34  ( .A(\i_iq_demod/filtre_I/current_state [2]), .B(\i_iq_demod/filtre_I/n6 ), .C(\i_iq_demod/filtre_I/n7 ), .Q(
        \i_iq_demod/filtre_I/n4 ) );
  DFEC1 \i_iq_demod/filtre_I/data_out_reg[0]  ( .D(
        \i_iq_demod/filtre_I/temp [9]), .E(\i_iq_demod/filtre_I/N123 ), .C(
        clk_i), .RN(resetn_i), .Q(demod_iq_ibb_o[0]) );
  DFEC1 \i_iq_demod/filtre_I/data_out_reg[1]  ( .D(
        \i_iq_demod/filtre_I/temp [10]), .E(\i_iq_demod/filtre_I/N123 ), .C(
        clk_i), .RN(resetn_i), .Q(demod_iq_ibb_o[1]) );
  DFEC1 \i_iq_demod/filtre_I/data_out_reg[2]  ( .D(
        \i_iq_demod/filtre_I/temp [11]), .E(\i_iq_demod/filtre_I/N123 ), .C(
        clk_i), .RN(resetn_i), .Q(demod_iq_ibb_o[2]) );
  DFEC1 \i_iq_demod/filtre_I/data_out_reg[3]  ( .D(
        \i_iq_demod/filtre_I/temp [12]), .E(\i_iq_demod/filtre_I/N123 ), .C(
        clk_i), .RN(resetn_i), .Q(demod_iq_ibb_o[3]) );
  DFEC1 \i_iq_demod/filtre_I/data_out_reg[4]  ( .D(
        \i_iq_demod/filtre_I/temp [13]), .E(\i_iq_demod/filtre_I/N123 ), .C(
        clk_i), .RN(resetn_i), .Q(demod_iq_ibb_o[4]) );
  DFC1 \i_iq_demod/filtre_I/out_valid_reg  ( .D(\i_iq_demod/filtre_I/N123 ), 
        .C(clk_i), .RN(resetn_i), .QN(n1412) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[13]  ( .D(\i_iq_demod/filtre_I/N28 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [13]) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[12]  ( .D(\i_iq_demod/filtre_I/N27 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [12]) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[11]  ( .D(\i_iq_demod/filtre_I/N26 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [11]), .QN(n249)
         );
  DFC1 \i_iq_demod/filtre_I/temp_reg[10]  ( .D(\i_iq_demod/filtre_I/N25 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [10]) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[9]  ( .D(\i_iq_demod/filtre_I/N24 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [9]), .QN(n250) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[8]  ( .D(\i_iq_demod/filtre_I/N23 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [8]) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[7]  ( .D(\i_iq_demod/filtre_I/N22 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [7]), .QN(n241) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[6]  ( .D(\i_iq_demod/filtre_I/N21 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [6]) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[5]  ( .D(\i_iq_demod/filtre_I/N20 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [5]), .QN(n242) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[4]  ( .D(\i_iq_demod/filtre_I/N19 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [4]) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[3]  ( .D(\i_iq_demod/filtre_I/N18 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [3]), .QN(n231) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[2]  ( .D(\i_iq_demod/filtre_I/N17 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [2]) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[1]  ( .D(\i_iq_demod/filtre_I/N16 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/temp [1]) );
  DFC1 \i_iq_demod/filtre_I/temp_reg[0]  ( .D(\i_iq_demod/filtre_I/N15 ), .C(
        clk_i), .RN(resetn_i), .QN(n228) );
  DFC1 \i_iq_demod/filtre_I/data_1_1_reg[4]  ( .D(
        \i_iq_demod/filtre_I/data_1_1_req [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_1_1 [4]) );
  DFC1 \i_iq_demod/filtre_I/data_1_1_reg[3]  ( .D(
        \i_iq_demod/filtre_I/data_1_1_req [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_1_1 [3]) );
  DFC1 \i_iq_demod/filtre_I/data_1_1_reg[2]  ( .D(
        \i_iq_demod/filtre_I/data_1_1_req [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_1_1 [2]) );
  DFC1 \i_iq_demod/filtre_I/data_2_1_reg[4]  ( .D(
        \i_iq_demod/filtre_I/data_2_1_req [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_2_1 [4]) );
  DFC1 \i_iq_demod/filtre_I/data_2_1_reg[3]  ( .D(
        \i_iq_demod/filtre_I/data_2_1_req [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_2_1 [3]) );
  DFC1 \i_iq_demod/filtre_I/data_2_1_reg[2]  ( .D(
        \i_iq_demod/filtre_I/data_2_1_req [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_2_1 [2]) );
  DFC1 \i_iq_demod/filtre_I/data_1_2_reg[4]  ( .D(
        \i_iq_demod/filtre_I/data_1_2_req [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_1_2 [4]) );
  DFC1 \i_iq_demod/filtre_I/data_1_2_reg[3]  ( .D(
        \i_iq_demod/filtre_I/data_1_2_req [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_1_2 [3]) );
  DFC1 \i_iq_demod/filtre_I/data_1_2_reg[2]  ( .D(
        \i_iq_demod/filtre_I/data_1_2_req [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_1_2 [2]) );
  DFC1 \i_iq_demod/filtre_I/data_2_2_reg[4]  ( .D(
        \i_iq_demod/filtre_I/data_2_2_req [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_2_2 [4]) );
  DFC1 \i_iq_demod/filtre_I/data_2_2_reg[3]  ( .D(
        \i_iq_demod/filtre_I/data_2_2_req [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_2_2 [3]) );
  DFC1 \i_iq_demod/filtre_I/data_2_2_reg[2]  ( .D(
        \i_iq_demod/filtre_I/data_2_2_req [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_2_2 [2]) );
  DFC1 \i_iq_demod/filtre_I/out_factor1_reg[8]  ( .D(
        \i_iq_demod/filtre_I/out_factor1_req [8]), .C(clk_i), .RN(resetn_i), 
        .QN(n212) );
  DFC1 \i_iq_demod/filtre_I/out_factor1_reg[7]  ( .D(
        \i_iq_demod/filtre_I/out_factor1_req [7]), .C(clk_i), .RN(resetn_i), 
        .QN(n208) );
  DFC1 \i_iq_demod/filtre_I/out_factor1_reg[6]  ( .D(
        \i_iq_demod/filtre_I/out_factor1_req [6]), .C(clk_i), .RN(resetn_i), 
        .Q(n1532), .QN(n156) );
  DFC1 \i_iq_demod/filtre_I/out_factor1_reg[5]  ( .D(
        \i_iq_demod/filtre_I/out_factor1_req [5]), .C(clk_i), .RN(resetn_i), 
        .QN(n142) );
  DFC1 \i_iq_demod/filtre_I/out_factor1_reg[0]  ( .D(
        \i_iq_demod/filtre_I/out_factor1_req [0]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_I/out_factor1 [0]), .QN(n146) );
  DFC1 \i_iq_demod/filtre_I/out_factor2_reg[8]  ( .D(
        \i_iq_demod/filtre_I/out_factor2_req [4]), .C(clk_i), .RN(resetn_i), 
        .QN(n175) );
  DFC1 \i_iq_demod/filtre_I/out_factor2_reg[7]  ( .D(
        \i_iq_demod/filtre_I/out_factor2_req [6]), .C(clk_i), .RN(resetn_i), 
        .QN(n171) );
  DFC1 \i_iq_demod/filtre_I/out_factor2_reg[6]  ( .D(
        \i_iq_demod/filtre_I/out_factor2_req [6]), .C(clk_i), .RN(resetn_i), 
        .QN(n169) );
  DFC1 \i_iq_demod/filtre_I/out_factor2_reg[5]  ( .D(
        \i_iq_demod/filtre_I/out_factor2_req [4]), .C(clk_i), .RN(resetn_i), 
        .QN(n139) );
  DFC1 \i_iq_demod/filtre_I/out_factor2_reg[0]  ( .D(
        \i_iq_demod/filtre_I/out_factor2_req [0]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_I/out_factor2 [0]), .QN(n143) );
  DFC3 \i_iq_demod/filtre_I/current_state_reg[1]  ( .D(
        \i_iq_demod/filtre_I/next_state [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/current_state [1]), .QN(\i_iq_demod/filtre_I/n6 )
         );
  DFC1 \i_iq_demod/filtre_I/current_state_reg[2]  ( .D(
        \i_iq_demod/filtre_I/sel [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/current_state [2]), .QN(\i_iq_demod/filtre_I/n2 )
         );
  DFC1 \i_iq_demod/filtre_I/current_state_reg[0]  ( .D(
        \i_iq_demod/filtre_I/next_state [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/current_state [0]) );
  NOR30 \i_iq_demod/gen_sin/U57  ( .A(\i_iq_demod/gen_sin/counter [0]), .B(
        \i_iq_demod/gen_sin/counter [1]), .C(\i_iq_demod/gen_sin/n22 ), .Q(
        \i_iq_demod/gen_sin/N106 ) );
  NOR20 \i_iq_demod/gen_sin/U56  ( .A(\i_iq_demod/gen_sin/N106 ), .B(
        \i_iq_demod/gen_sin/counter [0]), .Q(\i_iq_demod/gen_sin/N15 ) );
  NOR20 \i_iq_demod/gen_sin/U55  ( .A(\i_iq_demod/gen_sin/counter [1]), .B(
        \i_iq_demod/gen_sin/N106 ), .Q(\i_iq_demod/gen_sin/n21 ) );
  OAI210 \i_iq_demod/gen_sin/U54  ( .A(\i_iq_demod/gen_sin/n21 ), .B(
        \i_iq_demod/gen_sin/N15 ), .C(\i_iq_demod/gen_sin/counter [2]), .Q(
        \i_iq_demod/gen_sin/n20 ) );
  OAI310 \i_iq_demod/gen_sin/U53  ( .A(\i_iq_demod/gen_sin/n18 ), .B(
        \i_iq_demod/gen_sin/counter [2]), .C(\i_iq_demod/gen_sin/n19 ), .D(
        \i_iq_demod/gen_sin/n20 ), .Q(\i_iq_demod/gen_sin/N17 ) );
  CLKIN0 \i_iq_demod/gen_sin/U39  ( .A(\i_iq_demod/cosine_IN [1]), .Q(
        \i_iq_demod/gen_sin/n3 ) );
  CLKIN0 \i_iq_demod/gen_sin/U36  ( .A(\i_iq_demod/gen_sin/n6 ), .Q(
        \i_iq_demod/cosine_IN [0]) );
  OAI210 \i_iq_demod/gen_sin/U34  ( .A(\i_iq_demod/gen_sin/current_state [1]), 
        .B(\i_iq_demod/gen_sin/n1 ), .C(\i_iq_demod/gen_sin/n3 ), .Q(
        \i_iq_demod/gen_sin/next_state [1]) );
  NOR20 \i_iq_demod/gen_sin/U33  ( .A(\i_iq_demod/gen_sin/n2 ), .B(
        \i_iq_demod/gen_sin/n1 ), .Q(\i_iq_demod/sine_IN [1]) );
  CLKIN0 \i_iq_demod/gen_sin/U32  ( .A(\i_iq_demod/gen_sin/n1 ), .Q(
        \i_iq_demod/sine_IN [0]) );
  DFEC1 \i_iq_demod/gen_sin/current_state_reg[1]  ( .D(
        \i_iq_demod/gen_sin/next_state [1]), .E(\i_iq_demod/gen_sin/N106 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_iq_demod/gen_sin/current_state [1]), 
        .QN(\i_iq_demod/gen_sin/n2 ) );
  DFEC1 \i_iq_demod/gen_sin/current_state_reg[0]  ( .D(
        \i_iq_demod/gen_sin/next_state [0]), .E(\i_iq_demod/gen_sin/N106 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_iq_demod/gen_sin/current_state [0]) );
  DFC1 \i_iq_demod/gen_sin/counter_reg[2]  ( .D(\i_iq_demod/gen_sin/N17 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/gen_sin/counter [2]), .QN(
        \i_iq_demod/gen_sin/n22 ) );
  TFEC1 \i_iq_demod/gen_sin/counter_reg[1]  ( .T(
        \i_iq_demod/gen_sin/counter [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/gen_sin/counter [1]), .QN(\i_iq_demod/gen_sin/n18 ) );
  DFC3 \i_iq_demod/gen_sin/counter_reg[0]  ( .D(\i_iq_demod/gen_sin/N15 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/gen_sin/counter [0]), .QN(
        \i_iq_demod/gen_sin/n19 ) );
  NAND20 \i_cordic/S0/U43  ( .A(\i_cordic/S0/N9 ), .B(n1942), .Q(
        \i_cordic/S0/n37 ) );
  OAI210 \i_cordic/S0/U42  ( .A(n1942), .B(n276), .C(\i_cordic/S0/n37 ), .Q(
        \i_cordic/cor_x_s0[1][0] ) );
  CLKIN0 \i_cordic/S0/U41  ( .A(\i_cordic/S0/N4 ), .Q(\i_cordic/S0/n28 ) );
  CLKIN0 \i_cordic/S0/U38  ( .A(\i_cordic/S0/N5 ), .Q(\i_cordic/S0/n26 ) );
  NAND20 \i_cordic/S0/U37  ( .A(\i_cordic/S0/N11 ), .B(
        \i_cordic/cor_y_s0[0][5] ), .Q(\i_cordic/S0/n35 ) );
  CLKIN0 \i_cordic/S0/U35  ( .A(\i_cordic/S0/N6 ), .Q(\i_cordic/S0/n24 ) );
  NAND20 \i_cordic/S0/U34  ( .A(\i_cordic/S0/N12 ), .B(n1942), .Q(
        \i_cordic/S0/n34 ) );
  CLKIN0 \i_cordic/S0/U32  ( .A(\i_cordic/S0/N7 ), .Q(\i_cordic/S0/n22 ) );
  NAND20 \i_cordic/S0/U31  ( .A(\i_cordic/S0/N13 ), .B(n1942), .Q(
        \i_cordic/S0/n33 ) );
  OAI220 \i_cordic/S0/U25  ( .A(\i_cordic/S0/n39 ), .B(n276), .C(n1942), .D(
        n287), .Q(\i_cordic/cor_y_s0[1][0] ) );
  CLKIN0 \i_cordic/S0/U24  ( .A(\i_cordic/S0/N16 ), .Q(\i_cordic/S0/n29 ) );
  CLKIN0 \i_cordic/S0/U22  ( .A(\i_cordic/S0/N17 ), .Q(\i_cordic/S0/n27 ) );
  CLKIN0 \i_cordic/S0/U20  ( .A(\i_cordic/S0/N18 ), .Q(\i_cordic/S0/n25 ) );
  CLKIN0 \i_cordic/S0/U18  ( .A(\i_cordic/S0/N19 ), .Q(\i_cordic/S0/n23 ) );
  AOI220 \i_cordic/S1/U44  ( .A(n1942), .B(\i_cordic/S1/sub_50/B_not [5]), .C(
        n1942), .D(\i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/S1/n35 ) );
  CLKIN0 \i_cordic/S1/U43  ( .A(\i_cordic/S1/n35 ), .Q(
        \i_cordic/cor_w_s0[2][4] ) );
  AOI220 \i_cordic/S1/U42  ( .A(\i_cordic/S1/N38 ), .B(
        \i_cordic/S1/sub_50/B_not [5]), .C(\i_cordic/S1/N38 ), .D(
        \i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/S1/n34 ) );
  CLKIN0 \i_cordic/S1/U41  ( .A(\i_cordic/S1/n34 ), .Q(
        \i_cordic/cor_w_s0[2][5] ) );
  AOI220 \i_cordic/S2/U48  ( .A(\i_cordic/S2/N29 ), .B(n185), .C(n117), .D(
        \i_cordic/cor_y_s1[2][5] ), .Q(\i_cordic/S2/n37 ) );
  AOI220 \i_cordic/S2/U46  ( .A(\i_cordic/S2/N30 ), .B(n185), .C(
        \i_cordic/S2/N36 ), .D(\i_cordic/cor_y_s1[2][5] ), .Q(
        \i_cordic/S2/n36 ) );
  AOI220 \i_cordic/S2/U44  ( .A(\i_cordic/S2/N31 ), .B(n185), .C(
        \i_cordic/S2/N37 ), .D(\i_cordic/cor_y_s1[2][5] ), .Q(
        \i_cordic/S2/n35 ) );
  CLKIN0 \i_cordic/S2/U43  ( .A(\i_cordic/S2/n35 ), .Q(\i_cordic/S3/N37 ) );
  AOI220 \i_cordic/S2/U42  ( .A(\i_cordic/S2/N32 ), .B(n185), .C(
        \i_cordic/S2/N38 ), .D(\i_cordic/cor_y_s1[2][5] ), .Q(
        \i_cordic/S2/n34 ) );
  CLKIN0 \i_cordic/S2/U17  ( .A(\i_cordic/S2/n21 ), .Q(\i_cordic/S3/n30 ) );
  AOI220 \i_cordic/S3/U40  ( .A(\i_cordic/S3/N36 ), .B(\i_cordic/S2/n21 ), .C(
        \i_cordic/S3/N36 ), .D(\i_cordic/S3/n30 ), .Q(\i_cordic/S3/n28 ) );
  CLKIN0 \i_cordic/S3/U39  ( .A(\i_cordic/S3/n28 ), .Q(
        \i_cordic/cor_w_s1[4][3] ) );
  XNR20 \i_cdr/i_bit_recovery/U60  ( .A(\i_cdr/i_bit_recovery/phase_r [5]), 
        .B(\i_cdr/i_bit_recovery/phase_q [5]), .Q(\i_cdr/i_bit_recovery/n32 )
         );
  XOR20 \i_cdr/i_bit_recovery/U59  ( .A(\i_cdr/i_bit_recovery/phase_diff[5] ), 
        .B(\i_cdr/i_bit_recovery/phase_q [5]), .Q(\i_cdr/i_bit_recovery/n33 )
         );
  NAND20 \i_cdr/i_bit_recovery/U58  ( .A(\i_cdr/i_bit_recovery/n32 ), .B(
        \i_cdr/i_bit_recovery/n33 ), .Q(\i_cdr/i_bit_recovery/n31 ) );
  CLKIN0 \i_cdr/i_bit_recovery/U57  ( .A(\i_cdr/i_bit_recovery/n31 ), .Q(
        \i_cdr/i_bit_recovery/n25 ) );
  NOR30 \i_cdr/i_bit_recovery/U56  ( .A(\i_cdr/i_bit_recovery/phase_q [0]), 
        .B(\i_cdr/i_bit_recovery/phase_q [2]), .C(
        \i_cdr/i_bit_recovery/phase_q [1]), .Q(\i_cdr/i_bit_recovery/n27 ) );
  NOR30 \i_cdr/i_bit_recovery/U55  ( .A(\i_cdr/i_bit_recovery/phase_q [3]), 
        .B(\i_cdr/i_bit_recovery/phase_q [5]), .C(
        \i_cdr/i_bit_recovery/phase_q [4]), .Q(\i_cdr/i_bit_recovery/n28 ) );
  NOR30 \i_cdr/i_bit_recovery/U54  ( .A(\i_cdr/i_bit_recovery/phase_r [0]), 
        .B(\i_cdr/i_bit_recovery/phase_r [2]), .C(
        \i_cdr/i_bit_recovery/phase_r [1]), .Q(\i_cdr/i_bit_recovery/n29 ) );
  NOR30 \i_cdr/i_bit_recovery/U53  ( .A(\i_cdr/i_bit_recovery/phase_r [3]), 
        .B(\i_cdr/i_bit_recovery/phase_r [5]), .C(
        \i_cdr/i_bit_recovery/phase_r [4]), .Q(\i_cdr/i_bit_recovery/n30 ) );
  NAND40 \i_cdr/i_bit_recovery/U52  ( .A(\i_cdr/i_bit_recovery/n27 ), .B(
        \i_cdr/i_bit_recovery/n28 ), .C(\i_cdr/i_bit_recovery/n29 ), .D(
        \i_cdr/i_bit_recovery/n30 ), .Q(\i_cdr/i_bit_recovery/n26 ) );
  NOR20 \i_cdr/i_bit_recovery/U37  ( .A(\i_cdr/i_bit_recovery/curr_state [1]), 
        .B(\i_cdr/i_bit_recovery/n11 ), .Q(
        \i_cdr/i_bit_recovery/next_state [0]) );
  CLKIN0 \i_cdr/i_bit_recovery/U36  ( .A(cdr_valid_i), .Q(
        \i_cdr/i_bit_recovery/n9 ) );
  OAI220 \i_cdr/i_bit_recovery/U35  ( .A(\i_cdr/i_bit_recovery/n9 ), .B(
        \i_cdr/i_bit_recovery/n10 ), .C(\i_cdr/i_bit_recovery/n11 ), .D(
        \i_cdr/i_bit_recovery/n12 ), .Q(\i_cdr/i_bit_recovery/next_state [1])
         );
  INV2 \i_cdr/i_bit_recovery/U3  ( .A(\i_cdr/i_bit_recovery/phase_diff[5] ), 
        .Q(\i_cdr/i_bit_recovery/n8 ) );
  DLCQ3 \i_cdr/i_bit_recovery/data_bits_reg  ( .D(\i_cdr/i_bit_recovery/n8 ), 
        .GN(\i_cdr/i_bit_recovery/n25 ), .RN(\i_cdr/i_bit_recovery/n26 ), .Q(
        \i_cdr/data_w ) );
  DFEC1 \i_cdr/i_bit_recovery/phase_r_reg[0]  ( .D(
        \i_cdr/i_bit_recovery/phase_q [0]), .E(\i_cdr/i_bit_recovery/N91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_cdr/i_bit_recovery/phase_r [0]), .QN(
        n260) );
  DFEC1 \i_cdr/i_bit_recovery/phase_q_reg[0]  ( .D(cdr_phase_i[0]), .E(
        \i_cdr/i_bit_recovery/N91 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_cdr/i_bit_recovery/phase_q [0]) );
  DFEC1 \i_cdr/i_bit_recovery/phase_r_reg[1]  ( .D(
        \i_cdr/i_bit_recovery/phase_q [1]), .E(\i_cdr/i_bit_recovery/N91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_cdr/i_bit_recovery/phase_r [1]) );
  DFEC1 \i_cdr/i_bit_recovery/phase_q_reg[1]  ( .D(cdr_phase_i[1]), .E(
        \i_cdr/i_bit_recovery/N91 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_cdr/i_bit_recovery/phase_q [1]), .QN(n261) );
  DFEC1 \i_cdr/i_bit_recovery/phase_r_reg[2]  ( .D(
        \i_cdr/i_bit_recovery/phase_q [2]), .E(\i_cdr/i_bit_recovery/N91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_cdr/i_bit_recovery/phase_r [2]), .QN(
        n264) );
  DFEC1 \i_cdr/i_bit_recovery/phase_q_reg[2]  ( .D(cdr_phase_i[2]), .E(
        \i_cdr/i_bit_recovery/N91 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_cdr/i_bit_recovery/phase_q [2]) );
  DFEC1 \i_cdr/i_bit_recovery/phase_r_reg[3]  ( .D(
        \i_cdr/i_bit_recovery/phase_q [3]), .E(\i_cdr/i_bit_recovery/N91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_cdr/i_bit_recovery/phase_r [3]) );
  DFEC1 \i_cdr/i_bit_recovery/phase_q_reg[3]  ( .D(cdr_phase_i[3]), .E(
        \i_cdr/i_bit_recovery/N91 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_cdr/i_bit_recovery/phase_q [3]), .QN(n262) );
  DFEC1 \i_cdr/i_bit_recovery/phase_r_reg[4]  ( .D(
        \i_cdr/i_bit_recovery/phase_q [4]), .E(\i_cdr/i_bit_recovery/N91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_cdr/i_bit_recovery/phase_r [4]) );
  DFEC1 \i_cdr/i_bit_recovery/phase_q_reg[4]  ( .D(cdr_phase_i[4]), .E(
        \i_cdr/i_bit_recovery/N91 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_cdr/i_bit_recovery/phase_q [4]), .QN(n263) );
  DFEC1 \i_cdr/i_bit_recovery/phase_r_reg[5]  ( .D(
        \i_cdr/i_bit_recovery/phase_q [5]), .E(\i_cdr/i_bit_recovery/N91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_cdr/i_bit_recovery/phase_r [5]), .QN(
        n259) );
  DFEC1 \i_cdr/i_bit_recovery/phase_q_reg[5]  ( .D(cdr_phase_i[5]), .E(
        \i_cdr/i_bit_recovery/N91 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_cdr/i_bit_recovery/phase_q [5]) );
  DFC1 \i_cdr/i_bit_recovery/curr_state_reg[1]  ( .D(
        \i_cdr/i_bit_recovery/next_state [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_cdr/i_bit_recovery/curr_state [1]), .QN(\i_cdr/i_bit_recovery/n12 )
         );
  DFC3 \i_cdr/i_bit_recovery/curr_state_reg[0]  ( .D(
        \i_cdr/i_bit_recovery/next_state [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_cdr/i_bit_recovery/curr_state [0]), .QN(\i_cdr/i_bit_recovery/n14 )
         );
  NOR20 \i_cdr/i_cdr/U69  ( .A(\i_cdr/i_cdr/N145 ), .B(\i_cdr/i_cdr/count [0]), 
        .Q(\i_cdr/i_cdr/N153 ) );
  CLKIN0 \i_cdr/i_cdr/U68  ( .A(\i_cdr/i_cdr/N149 ), .Q(\i_cdr/i_cdr/n29 ) );
  NOR20 \i_cdr/i_cdr/U67  ( .A(\i_cdr/i_cdr/N145 ), .B(\i_cdr/i_cdr/n29 ), .Q(
        \i_cdr/i_cdr/N154 ) );
  CLKIN0 \i_cdr/i_cdr/U66  ( .A(\i_cdr/i_cdr/N150 ), .Q(\i_cdr/i_cdr/n28 ) );
  NOR20 \i_cdr/i_cdr/U65  ( .A(\i_cdr/i_cdr/N145 ), .B(\i_cdr/i_cdr/n28 ), .Q(
        \i_cdr/i_cdr/N155 ) );
  CLKIN0 \i_cdr/i_cdr/U64  ( .A(\i_cdr/i_cdr/N151 ), .Q(\i_cdr/i_cdr/n27 ) );
  NOR20 \i_cdr/i_cdr/U63  ( .A(\i_cdr/i_cdr/N145 ), .B(\i_cdr/i_cdr/n27 ), .Q(
        \i_cdr/i_cdr/N156 ) );
  NOR20 \i_cdr/i_cdr/U61  ( .A(\i_cdr/i_cdr/N145 ), .B(n246), .Q(
        \i_cdr/i_cdr/N157 ) );
  NOR30 \i_cdr/i_cdr/U42  ( .A(\i_cdr/i_cdr/count [0]), .B(
        \i_cdr/i_cdr/count [4]), .C(\i_cdr/i_cdr/count [1]), .Q(
        \i_cdr/i_cdr/n12 ) );
  AOI310 \i_cdr/i_cdr/U41  ( .A(\i_cdr/i_cdr/count [3]), .B(
        \i_cdr/i_cdr/count [2]), .C(\i_cdr/i_cdr/n12 ), .D(\i_cdr/i_cdr/N145 ), 
        .Q(\i_cdr/i_cdr/n11 ) );
  XOR20 \i_cdr/i_cdr/U40  ( .A(\i_cdr/i_cdr/q2 ), .B(\i_cdr/i_cdr/q1 ), .Q(
        \i_cdr/i_cdr/n9 ) );
  XNR20 \i_cdr/i_cdr/U38  ( .A(\i_cdr/i_cdr/q4 ), .B(\i_cdr/i_cdr/q2 ), .Q(
        \i_cdr/i_cdr/n4 ) );
  CLKIN0 \i_cdr/i_cdr/U37  ( .A(\i_cdr/i_cdr/n4 ), .Q(\i_cdr/i_cdr/n6 ) );
  NOR20 \i_cdr/i_cdr/U36  ( .A(\i_cdr/i_cdr/n5 ), .B(\i_cdr/i_cdr/n6 ), .Q(
        \i_cdr/i_cdr/next_state [0]) );
  NOR20 \i_cdr/i_cdr/U35  ( .A(\i_cdr/i_cdr/n4 ), .B(\i_cdr/i_cdr/n5 ), .Q(
        \i_cdr/i_cdr/next_state [1]) );
  INV2 \i_cdr/i_cdr/U3  ( .A(\i_cdr/i_cdr/n11 ), .Q(\i_cdr/i_cdr/n3 ) );
  DFC1 \i_cdr/i_cdr/data_en_o_reg  ( .D(\i_cdr/i_cdr/N160 ), .C(clk_i), .RN(
        resetn_i), .Q(cdr_valid_o), .QN(n186) );
  DFEC1 \i_cdr/i_cdr/data_o_reg  ( .D(\i_cdr/data_w ), .E(\i_cdr/i_cdr/N160 ), 
        .C(clk_i), .RN(resetn_i), .QN(n191) );
  DFC1 \i_cdr/i_cdr/data_en_w_q_reg  ( .D(\i_cdr/i_cdr/data_en_w ), .C(clk_i), 
        .RN(resetn_i), .QN(n121) );
  DFP1 \i_cdr/i_cdr/count_reg[3]  ( .D(\i_cdr/i_cdr/N156 ), .C(clk_i), .SN(
        resetn_i), .Q(\i_cdr/i_cdr/count [3]), .QN(n243) );
  DFC1 \i_cdr/i_cdr/count_reg[2]  ( .D(\i_cdr/i_cdr/N155 ), .C(clk_i), .RN(
        resetn_i), .Q(\i_cdr/i_cdr/count [2]) );
  DFC1 \i_cdr/i_cdr/count_reg[1]  ( .D(\i_cdr/i_cdr/N154 ), .C(clk_i), .RN(
        resetn_i), .Q(\i_cdr/i_cdr/count [1]), .QN(n116) );
  DFC1 \i_cdr/i_cdr/count_reg[0]  ( .D(\i_cdr/i_cdr/N153 ), .C(clk_i), .RN(
        resetn_i), .Q(\i_cdr/i_cdr/count [0]) );
  DFP1 \i_cdr/i_cdr/count_reg[4]  ( .D(\i_cdr/i_cdr/N157 ), .C(clk_i), .SN(
        resetn_i), .Q(\i_cdr/i_cdr/count [4]), .QN(n244) );
  DFC1 \i_cdr/i_cdr/curr_state_reg[1]  ( .D(\i_cdr/i_cdr/next_state [1]), .C(
        clk_i), .RN(resetn_i), .Q(\i_cdr/i_cdr/curr_state[1] ), .QN(
        \i_cdr/i_cdr/n8 ) );
  DFC3 \i_cdr/i_cdr/curr_state_reg[0]  ( .D(\i_cdr/i_cdr/next_state [0]), .C(
        clk_i), .RN(resetn_i), .QN(\i_cdr/i_cdr/n7 ) );
  DFC1 \i_cdr/i_cdr/q4_reg  ( .D(\i_cdr/i_cdr/q3 ), .C(\i_cdr/i_cdr/data_en_w ), .RN(resetn_i), .Q(\i_cdr/i_cdr/q4 ) );
  DFC1 \i_cdr/i_cdr/q3_reg  ( .D(\i_cdr/data_w ), .C(\i_cdr/i_cdr/N17 ), .RN(
        resetn_i), .Q(\i_cdr/i_cdr/q3 ) );
  DFC1 \i_cdr/i_cdr/q2_reg  ( .D(\i_cdr/i_cdr/q1 ), .C(\i_cdr/i_cdr/data_en_w ), .RN(resetn_i), .Q(\i_cdr/i_cdr/q2 ) );
  DFC1 \i_cdr/i_cdr/q1_reg  ( .D(\i_cdr/data_w ), .C(\i_cdr/i_cdr/data_en_w ), 
        .RN(resetn_i), .Q(\i_cdr/i_cdr/q1 ) );
  TFEP1 \i_cdr/i_cdr/data_en_w_reg  ( .T(\i_cdr/i_cdr/n3 ), .C(clk_i), .SN(
        resetn_i), .Q(\i_cdr/i_cdr/data_en_w ), .QN(\i_cdr/i_cdr/N17 ) );
  CLKIN0 \i_iq_demod/demod/validation/U36  ( .A(
        \i_iq_demod/demod/validation/n3 ), .Q(\i_iq_demod/filter_en ) );
  NOR20 \i_iq_demod/demod/validation/U34  ( .A(
        \i_iq_demod/demod/validation/current_state_valid [1]), .B(
        \i_iq_demod/demod/validation/n1 ), .Q(
        \i_iq_demod/demod/validation/next_state_valid [0]) );
  OAI210 \i_iq_demod/demod/validation/U33  ( .A(
        \i_iq_demod/demod/validation/n1 ), .B(\i_iq_demod/demod/validation/n2 ), .C(\i_iq_demod/demod/validation/n3 ), .Q(
        \i_iq_demod/demod/validation/next_state_valid [1]) );
  DFC1 \i_iq_demod/demod/validation/current_state_valid_reg[1]  ( .D(
        \i_iq_demod/demod/validation/next_state_valid [1]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/demod/validation/current_state_valid [1]), 
        .QN(\i_iq_demod/demod/validation/n2 ) );
  DFC3 \i_iq_demod/demod/validation/current_state_valid_reg[0]  ( .D(
        \i_iq_demod/demod/validation/next_state_valid [0]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/demod/validation/current_state_valid [0]), 
        .QN(\i_iq_demod/demod/validation/n5 ) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U44  ( .A(
        \i_iq_demod/filtre_I/shift_reg8 [0]), .B(
        \i_iq_demod/filtre_I/data_reg1/n7 ), .C(
        \i_iq_demod/filtre_I/shift_reg6 [0]), .D(
        \i_iq_demod/filtre_I/data_reg1/n8 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n33 ) );
  NAND20 \i_iq_demod/filtre_I/data_reg1/U42  ( .A(
        \i_iq_demod/filtre_I/shift_reg4 [0]), .B(
        \i_iq_demod/filtre_I/data_reg1/n6 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n34 ) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U39  ( .A(
        \i_iq_demod/filtre_I/shift_reg2 [0]), .B(
        \i_iq_demod/filtre_I/data_reg1/n4 ), .C(
        \i_iq_demod/filtre_I/shift_reg0 [0]), .D(
        \i_iq_demod/filtre_I/data_reg1/n5 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n35 ) );
  NAND30 \i_iq_demod/filtre_I/data_reg1/U38  ( .A(
        \i_iq_demod/filtre_I/data_reg1/n33 ), .B(
        \i_iq_demod/filtre_I/data_reg1/n34 ), .C(
        \i_iq_demod/filtre_I/data_reg1/n35 ), .Q(
        \i_iq_demod/filtre_I/data_1_1_req [0]) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U37  ( .A(
        \i_iq_demod/filtre_I/shift_reg8 [1]), .B(
        \i_iq_demod/filtre_I/data_reg1/n7 ), .C(
        \i_iq_demod/filtre_I/shift_reg6 [1]), .D(
        \i_iq_demod/filtre_I/data_reg1/n8 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n30 ) );
  NAND20 \i_iq_demod/filtre_I/data_reg1/U36  ( .A(
        \i_iq_demod/filtre_I/shift_reg4 [1]), .B(
        \i_iq_demod/filtre_I/data_reg1/n6 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n31 ) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U35  ( .A(
        \i_iq_demod/filtre_I/shift_reg2 [1]), .B(
        \i_iq_demod/filtre_I/data_reg1/n4 ), .C(
        \i_iq_demod/filtre_I/shift_reg0 [1]), .D(
        \i_iq_demod/filtre_I/data_reg1/n5 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n32 ) );
  NAND30 \i_iq_demod/filtre_I/data_reg1/U34  ( .A(
        \i_iq_demod/filtre_I/data_reg1/n30 ), .B(
        \i_iq_demod/filtre_I/data_reg1/n31 ), .C(
        \i_iq_demod/filtre_I/data_reg1/n32 ), .Q(
        \i_iq_demod/filtre_I/data_1_1_req [1]) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U33  ( .A(
        \i_iq_demod/filtre_I/shift_reg8 [2]), .B(
        \i_iq_demod/filtre_I/data_reg1/n7 ), .C(
        \i_iq_demod/filtre_I/shift_reg6 [2]), .D(
        \i_iq_demod/filtre_I/data_reg1/n8 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n27 ) );
  NAND20 \i_iq_demod/filtre_I/data_reg1/U32  ( .A(
        \i_iq_demod/filtre_I/shift_reg4 [2]), .B(
        \i_iq_demod/filtre_I/data_reg1/n6 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n28 ) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U31  ( .A(
        \i_iq_demod/filtre_I/shift_reg2 [2]), .B(
        \i_iq_demod/filtre_I/data_reg1/n4 ), .C(
        \i_iq_demod/filtre_I/shift_reg0 [2]), .D(
        \i_iq_demod/filtre_I/data_reg1/n5 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n29 ) );
  NAND30 \i_iq_demod/filtre_I/data_reg1/U30  ( .A(
        \i_iq_demod/filtre_I/data_reg1/n27 ), .B(
        \i_iq_demod/filtre_I/data_reg1/n28 ), .C(
        \i_iq_demod/filtre_I/data_reg1/n29 ), .Q(
        \i_iq_demod/filtre_I/data_1_1_req [2]) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U29  ( .A(
        \i_iq_demod/filtre_I/shift_reg8 [3]), .B(
        \i_iq_demod/filtre_I/data_reg1/n7 ), .C(
        \i_iq_demod/filtre_I/shift_reg6 [3]), .D(
        \i_iq_demod/filtre_I/data_reg1/n8 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n24 ) );
  NAND20 \i_iq_demod/filtre_I/data_reg1/U28  ( .A(
        \i_iq_demod/filtre_I/shift_reg4 [3]), .B(
        \i_iq_demod/filtre_I/data_reg1/n6 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n25 ) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U27  ( .A(
        \i_iq_demod/filtre_I/shift_reg2 [3]), .B(
        \i_iq_demod/filtre_I/data_reg1/n4 ), .C(
        \i_iq_demod/filtre_I/shift_reg0 [3]), .D(
        \i_iq_demod/filtre_I/data_reg1/n5 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n26 ) );
  NAND30 \i_iq_demod/filtre_I/data_reg1/U26  ( .A(
        \i_iq_demod/filtre_I/data_reg1/n24 ), .B(
        \i_iq_demod/filtre_I/data_reg1/n25 ), .C(
        \i_iq_demod/filtre_I/data_reg1/n26 ), .Q(
        \i_iq_demod/filtre_I/data_1_1_req [3]) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U25  ( .A(
        \i_iq_demod/filtre_I/shift_reg8 [4]), .B(
        \i_iq_demod/filtre_I/data_reg1/n7 ), .C(
        \i_iq_demod/filtre_I/shift_reg6 [4]), .D(
        \i_iq_demod/filtre_I/data_reg1/n8 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n21 ) );
  NAND20 \i_iq_demod/filtre_I/data_reg1/U24  ( .A(
        \i_iq_demod/filtre_I/shift_reg4 [4]), .B(
        \i_iq_demod/filtre_I/data_reg1/n6 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n22 ) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U23  ( .A(
        \i_iq_demod/filtre_I/shift_reg2 [4]), .B(
        \i_iq_demod/filtre_I/data_reg1/n4 ), .C(
        \i_iq_demod/filtre_I/shift_reg0 [4]), .D(
        \i_iq_demod/filtre_I/data_reg1/n5 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n23 ) );
  NAND30 \i_iq_demod/filtre_I/data_reg1/U22  ( .A(
        \i_iq_demod/filtre_I/data_reg1/n21 ), .B(
        \i_iq_demod/filtre_I/data_reg1/n22 ), .C(
        \i_iq_demod/filtre_I/data_reg1/n23 ), .Q(
        \i_iq_demod/filtre_I/data_1_1_req [4]) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U21  ( .A(
        \i_iq_demod/filtre_I/shift_reg9 [0]), .B(
        \i_iq_demod/filtre_I/data_reg1/n7 ), .C(
        \i_iq_demod/filtre_I/shift_reg7 [0]), .D(
        \i_iq_demod/filtre_I/data_reg1/n8 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n18 ) );
  NAND20 \i_iq_demod/filtre_I/data_reg1/U20  ( .A(
        \i_iq_demod/filtre_I/shift_reg5 [0]), .B(
        \i_iq_demod/filtre_I/data_reg1/n6 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n19 ) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U19  ( .A(
        \i_iq_demod/filtre_I/shift_reg3 [0]), .B(
        \i_iq_demod/filtre_I/data_reg1/n4 ), .C(
        \i_iq_demod/filtre_I/shift_reg1 [0]), .D(
        \i_iq_demod/filtre_I/data_reg1/n5 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n20 ) );
  NAND30 \i_iq_demod/filtre_I/data_reg1/U18  ( .A(
        \i_iq_demod/filtre_I/data_reg1/n18 ), .B(
        \i_iq_demod/filtre_I/data_reg1/n19 ), .C(
        \i_iq_demod/filtre_I/data_reg1/n20 ), .Q(
        \i_iq_demod/filtre_I/data_2_1_req [0]) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U17  ( .A(
        \i_iq_demod/filtre_I/shift_reg9 [1]), .B(
        \i_iq_demod/filtre_I/data_reg1/n7 ), .C(
        \i_iq_demod/filtre_I/shift_reg7 [1]), .D(
        \i_iq_demod/filtre_I/data_reg1/n8 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n15 ) );
  NAND20 \i_iq_demod/filtre_I/data_reg1/U16  ( .A(
        \i_iq_demod/filtre_I/shift_reg5 [1]), .B(
        \i_iq_demod/filtre_I/data_reg1/n6 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n16 ) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U15  ( .A(
        \i_iq_demod/filtre_I/shift_reg3 [1]), .B(
        \i_iq_demod/filtre_I/data_reg1/n4 ), .C(
        \i_iq_demod/filtre_I/shift_reg1 [1]), .D(
        \i_iq_demod/filtre_I/data_reg1/n5 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n17 ) );
  NAND30 \i_iq_demod/filtre_I/data_reg1/U14  ( .A(
        \i_iq_demod/filtre_I/data_reg1/n15 ), .B(
        \i_iq_demod/filtre_I/data_reg1/n16 ), .C(
        \i_iq_demod/filtre_I/data_reg1/n17 ), .Q(
        \i_iq_demod/filtre_I/data_2_1_req [1]) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U13  ( .A(
        \i_iq_demod/filtre_I/shift_reg9 [2]), .B(
        \i_iq_demod/filtre_I/data_reg1/n7 ), .C(
        \i_iq_demod/filtre_I/shift_reg7 [2]), .D(
        \i_iq_demod/filtre_I/data_reg1/n8 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n12 ) );
  NAND20 \i_iq_demod/filtre_I/data_reg1/U12  ( .A(
        \i_iq_demod/filtre_I/shift_reg5 [2]), .B(
        \i_iq_demod/filtre_I/data_reg1/n6 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n13 ) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U11  ( .A(
        \i_iq_demod/filtre_I/shift_reg3 [2]), .B(
        \i_iq_demod/filtre_I/data_reg1/n4 ), .C(
        \i_iq_demod/filtre_I/shift_reg1 [2]), .D(
        \i_iq_demod/filtre_I/data_reg1/n5 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n14 ) );
  NAND30 \i_iq_demod/filtre_I/data_reg1/U10  ( .A(
        \i_iq_demod/filtre_I/data_reg1/n12 ), .B(
        \i_iq_demod/filtre_I/data_reg1/n13 ), .C(
        \i_iq_demod/filtre_I/data_reg1/n14 ), .Q(
        \i_iq_demod/filtre_I/data_2_1_req [2]) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U9  ( .A(
        \i_iq_demod/filtre_I/shift_reg9 [3]), .B(
        \i_iq_demod/filtre_I/data_reg1/n7 ), .C(
        \i_iq_demod/filtre_I/shift_reg7 [3]), .D(
        \i_iq_demod/filtre_I/data_reg1/n8 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n9 ) );
  NAND20 \i_iq_demod/filtre_I/data_reg1/U8  ( .A(
        \i_iq_demod/filtre_I/shift_reg5 [3]), .B(
        \i_iq_demod/filtre_I/data_reg1/n6 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n10 ) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U7  ( .A(
        \i_iq_demod/filtre_I/shift_reg3 [3]), .B(
        \i_iq_demod/filtre_I/data_reg1/n4 ), .C(
        \i_iq_demod/filtre_I/shift_reg1 [3]), .D(
        \i_iq_demod/filtre_I/data_reg1/n5 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n11 ) );
  NAND30 \i_iq_demod/filtre_I/data_reg1/U6  ( .A(
        \i_iq_demod/filtre_I/data_reg1/n9 ), .B(
        \i_iq_demod/filtre_I/data_reg1/n10 ), .C(
        \i_iq_demod/filtre_I/data_reg1/n11 ), .Q(
        \i_iq_demod/filtre_I/data_2_1_req [3]) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U5  ( .A(
        \i_iq_demod/filtre_I/shift_reg9 [4]), .B(
        \i_iq_demod/filtre_I/data_reg1/n7 ), .C(
        \i_iq_demod/filtre_I/shift_reg7 [4]), .D(
        \i_iq_demod/filtre_I/data_reg1/n8 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n1 ) );
  NAND20 \i_iq_demod/filtre_I/data_reg1/U4  ( .A(
        \i_iq_demod/filtre_I/shift_reg5 [4]), .B(
        \i_iq_demod/filtre_I/data_reg1/n6 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n2 ) );
  AOI220 \i_iq_demod/filtre_I/data_reg1/U3  ( .A(
        \i_iq_demod/filtre_I/shift_reg3 [4]), .B(
        \i_iq_demod/filtre_I/data_reg1/n4 ), .C(
        \i_iq_demod/filtre_I/shift_reg1 [4]), .D(
        \i_iq_demod/filtre_I/data_reg1/n5 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n3 ) );
  NAND30 \i_iq_demod/filtre_I/data_reg1/U2  ( .A(
        \i_iq_demod/filtre_I/data_reg1/n1 ), .B(
        \i_iq_demod/filtre_I/data_reg1/n2 ), .C(
        \i_iq_demod/filtre_I/data_reg1/n3 ), .Q(
        \i_iq_demod/filtre_I/data_2_1_req [4]) );
  NOR30 \i_iq_demod/filtre_I/factor/U75  ( .A(\i_iq_demod/filtre_I/sel [0]), 
        .B(n1943), .C(\i_iq_demod/filtre_I/n9 ), .Q(
        \i_iq_demod/filtre_I/factor/n6 ) );
  NAND20 \i_iq_demod/filtre_I/shift_r/U9  ( .A(
        \i_iq_demod/filtre_I/shift_count [0]), .B(
        \i_iq_demod/filtre_I/shift_count [1]), .Q(
        \i_iq_demod/filtre_I/shift_r/n5 ) );
  XNR20 \i_iq_demod/filtre_I/shift_r/U7  ( .A(\i_iq_demod/filtre_I/shift_r/n1 ), .B(\i_iq_demod/filtre_I/shift_count [0]), .Q(
        \i_iq_demod/filtre_I/shift_r/N9 ) );
  AOI210 \i_iq_demod/filtre_I/shift_r/U6  ( .A(
        \i_iq_demod/filtre_I/shift_r/n5 ), .B(\i_iq_demod/demod/validation/n3 ), .C(\i_iq_demod/filtre_I/shift_r/N9 ), .Q(\i_iq_demod/filtre_I/shift_r/n6 )
         );
  CLKIN0 \i_iq_demod/filtre_I/shift_r/U5  ( .A(
        \i_iq_demod/filtre_I/shift_r/n5 ), .Q(\i_iq_demod/filtre_I/shift_r/n2 ) );
  NOR40 \i_iq_demod/filtre_I/shift_r/U4  ( .A(\i_iq_demod/filtre_I/shift_r/n2 ), .B(\i_iq_demod/filtre_I/shift_r/N9 ), .C(\i_iq_demod/filtre_I/shift_r/n3 ), 
        .D(\i_iq_demod/demod/validation/n3 ), .Q(
        \i_iq_demod/filtre_I/shift_r/N3 ) );
  AOI310 \i_iq_demod/filtre_I/shift_r/U3  ( .A(
        \i_iq_demod/filtre_I/shift_count [2]), .B(
        \i_iq_demod/filtre_I/shift_r/n1 ), .C(\i_iq_demod/filter_en ), .D(
        \i_iq_demod/filtre_I/shift_count [0]), .Q(
        \i_iq_demod/filtre_I/shift_r/N8 ) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out19_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg18 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg19 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out18_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg17 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg18 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out17_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg16 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg17 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out16_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg15 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg16 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out15_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg14 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg15 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out14_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg13 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg14 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out13_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg12 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg13 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out12_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg11 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg12 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out11_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg10 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg11 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out10_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg9 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg10 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out9_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg8 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg9 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out8_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg7 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg8 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out7_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg6 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg7 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out6_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg5 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg6 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out5_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg4 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg5 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out4_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg3 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg4 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out3_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg2 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg3 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out2_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg1 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg2 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out1_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_reg0 [0]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg1 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out0_reg[0]  ( .D(
        \i_iq_demod/I_BB_IN [0]), .E(n268), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/shift_reg0 [0]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out19_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg18 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg19 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out18_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg17 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg18 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out17_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg16 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg17 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out16_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg15 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg16 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out15_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg14 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg15 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out14_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg13 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg14 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out13_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg12 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg13 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out12_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg11 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg12 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out11_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg10 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg11 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out10_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg9 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg10 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out9_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg8 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg9 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out8_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg7 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg8 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out7_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg6 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg7 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out6_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg5 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg6 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out5_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg4 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg5 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out4_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg3 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg4 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out3_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg2 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg3 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out2_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg1 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg2 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out1_reg[1]  ( .D(
        \i_iq_demod/filtre_I/shift_reg0 [1]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg1 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out0_reg[1]  ( .D(
        \i_iq_demod/I_BB_IN [1]), .E(n268), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/shift_reg0 [1]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out19_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg18 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg19 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out18_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg17 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg18 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out17_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg16 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg17 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out16_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg15 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg16 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out15_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg14 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg15 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out14_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg13 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg14 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out13_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg12 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg13 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out12_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg11 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg12 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out11_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg10 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg11 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out10_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg9 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg10 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out9_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg8 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg9 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out8_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg7 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg8 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out7_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg6 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg7 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out6_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg5 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg6 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out5_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg4 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg5 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out4_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg3 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg4 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out3_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg2 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg3 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out2_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg1 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg2 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out1_reg[2]  ( .D(
        \i_iq_demod/filtre_I/shift_reg0 [2]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg1 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out0_reg[2]  ( .D(
        \i_iq_demod/I_BB_IN [2]), .E(n268), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/shift_reg0 [2]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out19_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg18 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg19 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out18_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg17 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg18 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out17_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg16 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg17 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out16_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg15 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg16 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out15_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg14 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg15 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out14_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg13 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg14 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out13_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg12 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg13 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out12_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg11 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg12 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out11_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg10 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg11 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out10_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg9 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg10 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out9_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg8 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg9 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out8_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg7 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg8 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out7_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg6 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg7 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out6_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg5 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg6 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out5_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg4 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg5 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out4_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg3 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg4 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out3_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg2 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg3 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out2_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg1 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg2 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out1_reg[3]  ( .D(
        \i_iq_demod/filtre_I/shift_reg0 [3]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg1 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out0_reg[3]  ( .D(
        \i_iq_demod/I_BB_IN [3]), .E(n268), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/shift_reg0 [3]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out19_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg18 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg19 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out18_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg17 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg18 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out17_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg16 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg17 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out16_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg15 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg16 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out15_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg14 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg15 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out14_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg13 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg14 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out13_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg12 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg13 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out12_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg11 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg12 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out11_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg10 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg11 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out10_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg9 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg10 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out9_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg8 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg9 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out8_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg7 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg8 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out7_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg6 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg7 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out6_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg5 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg6 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out5_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg4 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg5 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out4_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg3 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg4 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out3_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg2 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg3 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out2_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg1 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg2 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out1_reg[4]  ( .D(
        \i_iq_demod/filtre_I/shift_reg0 [4]), .E(n268), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/shift_reg1 [4]) );
  DFEC1 \i_iq_demod/filtre_I/shift_r/data_out0_reg[4]  ( .D(
        \i_iq_demod/I_BB_IN [4]), .E(n268), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/shift_reg0 [4]) );
  JKC1 \i_iq_demod/filtre_I/shift_r/cpt_shift_reg[2]  ( .J(
        \i_iq_demod/filtre_I/shift_r/n2 ), .K(\i_iq_demod/filtre_I/shift_r/n6 ), .C(clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_I/shift_count [2]), .QN(
        \i_iq_demod/filtre_I/shift_r/n3 ) );
  TFEC3 \i_iq_demod/filtre_I/shift_r/cpt_shift_reg[1]  ( .T(
        \i_iq_demod/filtre_I/shift_count [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/shift_count [1]), .QN(
        \i_iq_demod/filtre_I/shift_r/n1 ) );
  DFC1 \i_iq_demod/filtre_I/shift_r/cpt_shift_reg[0]  ( .D(
        \i_iq_demod/filtre_I/shift_r/N8 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/shift_count [0]) );
  XNR20 \i_iq_demod/filtre_I/temp_adder/U75  ( .A(n228), .B(
        \i_iq_demod/filtre_I/tot [0]), .Q(\i_iq_demod/filtre_I/n_temp [0]) );
  CLKIN0 \i_iq_demod/filtre_I/temp_adder/U74  ( .A(
        \i_iq_demod/filtre_I/tot [9]), .Q(\i_iq_demod/filtre_I/temp_adder/n45 ) );
  CLKIN0 \i_iq_demod/filtre_I/temp_adder/U72  ( .A(
        \i_iq_demod/filtre_I/tot [7]), .Q(\i_iq_demod/filtre_I/temp_adder/n48 ) );
  CLKIN0 \i_iq_demod/filtre_I/temp_adder/U70  ( .A(
        \i_iq_demod/filtre_I/tot [5]), .Q(\i_iq_demod/filtre_I/temp_adder/n51 ) );
  CLKIN0 \i_iq_demod/filtre_I/temp_adder/U68  ( .A(
        \i_iq_demod/filtre_I/tot [3]), .Q(\i_iq_demod/filtre_I/temp_adder/n54 ) );
  CLKIN0 \i_iq_demod/filtre_I/temp_adder/U66  ( .A(
        \i_iq_demod/filtre_I/tot [0]), .Q(\i_iq_demod/filtre_I/temp_adder/n20 ) );
  XNR20 \i_iq_demod/filtre_I/temp_adder/U65  ( .A(\i_iq_demod/filtre_I/tot [1]), .B(\i_iq_demod/filtre_I/temp [1]), .Q(\i_iq_demod/filtre_I/temp_adder/n17 )
         );
  NAND20 \i_iq_demod/filtre_I/temp_adder/U64  ( .A(
        \i_iq_demod/filtre_I/temp [1]), .B(\i_iq_demod/filtre_I/tot [1]), .Q(
        \i_iq_demod/filtre_I/temp_adder/n57 ) );
  OAI310 \i_iq_demod/filtre_I/temp_adder/U63  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n20 ), .B(
        \i_iq_demod/filtre_I/temp_adder/n17 ), .C(n228), .D(
        \i_iq_demod/filtre_I/temp_adder/n57 ), .Q(
        \i_iq_demod/filtre_I/temp_adder/n15 ) );
  XNR20 \i_iq_demod/filtre_I/temp_adder/U59  ( .A(\i_iq_demod/filtre_I/tot [3]), .B(\i_iq_demod/filtre_I/temp [3]), .Q(\i_iq_demod/filtre_I/temp_adder/n14 )
         );
  OAI220 \i_iq_demod/filtre_I/temp_adder/U58  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n54 ), .B(n231), .C(
        \i_iq_demod/filtre_I/temp_adder/n13 ), .D(
        \i_iq_demod/filtre_I/temp_adder/n14 ), .Q(
        \i_iq_demod/filtre_I/temp_adder/n11 ) );
  XNR20 \i_iq_demod/filtre_I/temp_adder/U54  ( .A(\i_iq_demod/filtre_I/tot [5]), .B(\i_iq_demod/filtre_I/temp [5]), .Q(\i_iq_demod/filtre_I/temp_adder/n10 )
         );
  OAI220 \i_iq_demod/filtre_I/temp_adder/U53  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n51 ), .B(n242), .C(
        \i_iq_demod/filtre_I/temp_adder/n9 ), .D(
        \i_iq_demod/filtre_I/temp_adder/n10 ), .Q(
        \i_iq_demod/filtre_I/temp_adder/n7 ) );
  XNR20 \i_iq_demod/filtre_I/temp_adder/U49  ( .A(\i_iq_demod/filtre_I/tot [7]), .B(\i_iq_demod/filtre_I/temp [7]), .Q(\i_iq_demod/filtre_I/temp_adder/n6 )
         );
  OAI220 \i_iq_demod/filtre_I/temp_adder/U48  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n48 ), .B(n241), .C(
        \i_iq_demod/filtre_I/temp_adder/n5 ), .D(
        \i_iq_demod/filtre_I/temp_adder/n6 ), .Q(
        \i_iq_demod/filtre_I/temp_adder/n3 ) );
  XNR20 \i_iq_demod/filtre_I/temp_adder/U44  ( .A(\i_iq_demod/filtre_I/tot [9]), .B(\i_iq_demod/filtre_I/temp [9]), .Q(\i_iq_demod/filtre_I/temp_adder/n2 )
         );
  OAI220 \i_iq_demod/filtre_I/temp_adder/U43  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n45 ), .B(n250), .C(
        \i_iq_demod/filtre_I/temp_adder/n1 ), .D(
        \i_iq_demod/filtre_I/temp_adder/n2 ), .Q(
        \i_iq_demod/filtre_I/temp_adder/n42 ) );
  XNR20 \i_iq_demod/filtre_I/temp_adder/U38  ( .A(
        \i_iq_demod/filtre_I/tot [11]), .B(\i_iq_demod/filtre_I/temp [11]), 
        .Q(\i_iq_demod/filtre_I/temp_adder/n41 ) );
  XOR20 \i_iq_demod/filtre_I/temp_adder/U37  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n40 ), .B(
        \i_iq_demod/filtre_I/temp_adder/n41 ), .Q(
        \i_iq_demod/filtre_I/n_temp [11]) );
  CLKIN0 \i_iq_demod/filtre_I/temp_adder/U36  ( .A(
        \i_iq_demod/filtre_I/tot [11]), .Q(
        \i_iq_demod/filtre_I/temp_adder/n38 ) );
  OAI220 \i_iq_demod/filtre_I/temp_adder/U34  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n38 ), .B(n249), .C(
        \i_iq_demod/filtre_I/temp_adder/n40 ), .D(
        \i_iq_demod/filtre_I/temp_adder/n41 ), .Q(
        \i_iq_demod/filtre_I/temp_adder/n35 ) );
  NOR20 \i_iq_demod/filtre_I/temp_adder/U11  ( .A(n228), .B(
        \i_iq_demod/filtre_I/temp_adder/n20 ), .Q(
        \i_iq_demod/filtre_I/temp_adder/n18 ) );
  XNR20 \i_iq_demod/filtre_I/temp_adder/U10  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n17 ), .B(
        \i_iq_demod/filtre_I/temp_adder/n18 ), .Q(
        \i_iq_demod/filtre_I/n_temp [1]) );
  XOR20 \i_iq_demod/filtre_I/temp_adder/U8  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n13 ), .B(
        \i_iq_demod/filtre_I/temp_adder/n14 ), .Q(
        \i_iq_demod/filtre_I/n_temp [3]) );
  XOR20 \i_iq_demod/filtre_I/temp_adder/U6  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n9 ), .B(
        \i_iq_demod/filtre_I/temp_adder/n10 ), .Q(
        \i_iq_demod/filtre_I/n_temp [5]) );
  XOR20 \i_iq_demod/filtre_I/temp_adder/U4  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n5 ), .B(
        \i_iq_demod/filtre_I/temp_adder/n6 ), .Q(
        \i_iq_demod/filtre_I/n_temp [7]) );
  XOR20 \i_iq_demod/filtre_I/temp_adder/U2  ( .A(
        \i_iq_demod/filtre_I/temp_adder/n1 ), .B(
        \i_iq_demod/filtre_I/temp_adder/n2 ), .Q(
        \i_iq_demod/filtre_I/n_temp [9]) );
  XOR20 \i_iq_demod/filtre_I/sum1_adder/U10  ( .A(
        \i_iq_demod/filtre_I/data_2_1 [3]), .B(
        \i_iq_demod/filtre_I/data_1_1 [3]), .Q(
        \i_iq_demod/filtre_I/sum1_adder/n6 ) );
  CLKIN0 \i_iq_demod/filtre_I/sum1_adder/U8  ( .A(
        \i_iq_demod/filtre_I/sum1_adder/n7 ), .Q(
        \i_iq_demod/filtre_I/sum1_adder/n5 ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U107  ( .A(n142), .B(n138), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[5] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U105  ( .A(n156), .B(n138), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[6] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U103  ( .A(n208), .B(n138), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[1][6] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U101  ( .A(n138), .B(n212), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[1][7] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U97  ( .A(n201), .B(n174), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[2] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U95  ( .A(n154), .B(n174), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[4] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U92  ( .A(n208), .B(n174), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[7] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U91  ( .A(n174), .B(n212), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[9] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U89  ( .A(n146), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[0] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U87  ( .A(n201), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[2] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U86  ( .A(n130), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[3] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U85  ( .A(n154), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[4] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U82  ( .A(n208), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[7] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U81  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .B(n212), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[9] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U78  ( .A(n202), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[1] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U77  ( .A(n201), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[2] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U76  ( .A(n130), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[3] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U75  ( .A(n154), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[4] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U72  ( .A(n208), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[7] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U68  ( .A(n202), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[1] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U67  ( .A(n201), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[2] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U65  ( .A(n154), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[4] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U63  ( .A(n156), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[6] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U58  ( .A(n202), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[1] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U57  ( .A(n201), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[2] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U56  ( .A(n130), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[3] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U55  ( .A(n154), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[4] ) );
  NAND20 \i_iq_demod/filtre_I/mult1_multiplier/U48  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/A_pipe [1]), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/B_pipe ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/n20 ) );
  NAND20 \i_iq_demod/filtre_I/mult1_multiplier/U46  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/A_pipe [2]), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/B_pipe ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/n19 ) );
  CLKIN0 \i_iq_demod/filtre_I/mult1_multiplier/U45  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/n19 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[2] ) );
  NAND20 \i_iq_demod/filtre_I/mult1_multiplier/U44  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/A_pipe [3]), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/B_pipe ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/n18 ) );
  CLKIN0 \i_iq_demod/filtre_I/mult1_multiplier/U43  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/n18 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[3] ) );
  NAND20 \i_iq_demod/filtre_I/mult1_multiplier/U42  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/A_pipe [4]), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/B_pipe ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/n17 ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U25  ( .A(n156), .B(n1709), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[6] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U24  ( .A(n208), .B(net42978), 
        .Q(\i_iq_demod/filtre_I/mult1_multiplier/_3_net_[7] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U23  ( .A(net42978), .B(n212), 
        .Q(\i_iq_demod/filtre_I/mult1_multiplier/_3_net_[9] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U16  ( .A(n142), .B(n166), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[5] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U14  ( .A(n208), .B(n166), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[7] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U8  ( .A(n168), .B(n130), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[3] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U6  ( .A(n168), .B(n142), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[5] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U5  ( .A(n168), .B(n156), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[6] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U4  ( .A(n168), .B(n208), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[7] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U3  ( .A(n168), .B(n212), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[9] ) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/B_pipe_reg  ( .D(
        \i_iq_demod/filtre_I/_15_net_[8] ), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/B_pipe ) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/A_pipe_reg[0]  ( .D(
        \i_iq_demod/filtre_I/out_factor1 [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/A_pipe [0]) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/A_pipe_reg[1]  ( .D(
        \i_iq_demod/filtre_I/out_factor1 [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/A_pipe [1]) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/A_pipe_reg[2]  ( .D(
        \i_iq_demod/filtre_I/out_factor1 [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/A_pipe [2]) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/A_pipe_reg[3]  ( .D(
        \i_iq_demod/filtre_I/out_factor1 [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/A_pipe [3]) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/A_pipe_reg[4]  ( .D(
        \i_iq_demod/filtre_I/out_factor1 [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/A_pipe [4]) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/register_pipe_reg[9][0]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/register[9][0] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][0] ), .QN(n214)
         );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/register_pipe_reg[9][1]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/register[9][1] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][1] ) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/register_pipe_reg[9][2]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/register[9][2] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][2] ) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/register_pipe_reg[9][3]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/register[9][3] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][3] ), .QN(n219)
         );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/register_pipe_reg[9][4]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/register[9][4] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][4] ) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/S_reg[0]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[0] ), .C(clk_i), .RN(
        resetn_i), .QN(n158) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/S_reg[1]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [1]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult1 [1]) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/S_reg[2]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [2]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult1 [2]) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/S_reg[3]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [3]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult1 [3]), .QN(n184) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/S_reg[4]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [4]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult1 [4]) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/S_reg[5]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [5]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult1 [5]), .QN(n190) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/S_reg[6]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [6]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult1 [6]) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/S_reg[7]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [7]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult1 [7]), .QN(n189) );
  DFC1 \i_iq_demod/filtre_I/mult1_multiplier/S_reg[8]  ( .D(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [8]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult1 [8]) );
  XNR20 \i_iq_demod/filtre_I/tot_adder/U66  ( .A(n158), .B(
        \i_iq_demod/filtre_I/mult2 [0]), .Q(\i_iq_demod/filtre_I/tot [0]) );
  CLKIN0 \i_iq_demod/filtre_I/tot_adder/U65  ( .A(
        \i_iq_demod/filtre_I/mult2 [9]), .Q(
        \i_iq_demod/filtre_I/tot_adder/n38 ) );
  CLKIN0 \i_iq_demod/filtre_I/tot_adder/U64  ( .A(
        \i_iq_demod/filtre_I/mult1 [9]), .Q(
        \i_iq_demod/filtre_I/tot_adder/n39 ) );
  XNR20 \i_iq_demod/filtre_I/tot_adder/U56  ( .A(
        \i_iq_demod/filtre_I/mult2 [1]), .B(\i_iq_demod/filtre_I/mult1 [1]), 
        .Q(\i_iq_demod/filtre_I/tot_adder/n17 ) );
  NAND20 \i_iq_demod/filtre_I/tot_adder/U55  ( .A(
        \i_iq_demod/filtre_I/mult1 [1]), .B(\i_iq_demod/filtre_I/mult2 [1]), 
        .Q(\i_iq_demod/filtre_I/tot_adder/n50 ) );
  OAI310 \i_iq_demod/filtre_I/tot_adder/U54  ( .A(n181), .B(
        \i_iq_demod/filtre_I/tot_adder/n17 ), .C(n158), .D(
        \i_iq_demod/filtre_I/tot_adder/n50 ), .Q(
        \i_iq_demod/filtre_I/tot_adder/n15 ) );
  XNR20 \i_iq_demod/filtre_I/tot_adder/U50  ( .A(
        \i_iq_demod/filtre_I/mult2 [3]), .B(\i_iq_demod/filtre_I/mult1 [3]), 
        .Q(\i_iq_demod/filtre_I/tot_adder/n14 ) );
  OAI220 \i_iq_demod/filtre_I/tot_adder/U49  ( .A(n224), .B(n184), .C(
        \i_iq_demod/filtre_I/tot_adder/n13 ), .D(
        \i_iq_demod/filtre_I/tot_adder/n14 ), .Q(
        \i_iq_demod/filtre_I/tot_adder/n11 ) );
  XNR20 \i_iq_demod/filtre_I/tot_adder/U45  ( .A(
        \i_iq_demod/filtre_I/mult2 [5]), .B(\i_iq_demod/filtre_I/mult1 [5]), 
        .Q(\i_iq_demod/filtre_I/tot_adder/n10 ) );
  OAI220 \i_iq_demod/filtre_I/tot_adder/U44  ( .A(n235), .B(n190), .C(
        \i_iq_demod/filtre_I/tot_adder/n9 ), .D(
        \i_iq_demod/filtre_I/tot_adder/n10 ), .Q(
        \i_iq_demod/filtre_I/tot_adder/n7 ) );
  XNR20 \i_iq_demod/filtre_I/tot_adder/U40  ( .A(
        \i_iq_demod/filtre_I/mult2 [7]), .B(\i_iq_demod/filtre_I/mult1 [7]), 
        .Q(\i_iq_demod/filtre_I/tot_adder/n6 ) );
  OAI220 \i_iq_demod/filtre_I/tot_adder/U39  ( .A(n234), .B(n189), .C(
        \i_iq_demod/filtre_I/tot_adder/n5 ), .D(
        \i_iq_demod/filtre_I/tot_adder/n6 ), .Q(
        \i_iq_demod/filtre_I/tot_adder/n3 ) );
  XNR20 \i_iq_demod/filtre_I/tot_adder/U35  ( .A(
        \i_iq_demod/filtre_I/mult2 [9]), .B(\i_iq_demod/filtre_I/mult1 [9]), 
        .Q(\i_iq_demod/filtre_I/tot_adder/n2 ) );
  OAI220 \i_iq_demod/filtre_I/tot_adder/U34  ( .A(
        \i_iq_demod/filtre_I/tot_adder/n38 ), .B(
        \i_iq_demod/filtre_I/tot_adder/n39 ), .C(
        \i_iq_demod/filtre_I/tot_adder/n1 ), .D(
        \i_iq_demod/filtre_I/tot_adder/n2 ), .Q(
        \i_iq_demod/filtre_I/tot_adder/n35 ) );
  XNR20 \i_iq_demod/filtre_I/tot_adder/U29  ( .A(
        \i_iq_demod/filtre_I/mult2 [11]), .B(\i_iq_demod/filtre_I/mult1 [11]), 
        .Q(\i_iq_demod/filtre_I/tot_adder/n34 ) );
  XOR20 \i_iq_demod/filtre_I/tot_adder/U28  ( .A(
        \i_iq_demod/filtre_I/tot_adder/n33 ), .B(
        \i_iq_demod/filtre_I/tot_adder/n34 ), .Q(\i_iq_demod/filtre_I/tot [11]) );
  CLKIN0 \i_iq_demod/filtre_I/tot_adder/U27  ( .A(
        \i_iq_demod/filtre_I/mult2 [11]), .Q(
        \i_iq_demod/filtre_I/tot_adder/n31 ) );
  CLKIN0 \i_iq_demod/filtre_I/tot_adder/U26  ( .A(
        \i_iq_demod/filtre_I/mult1 [11]), .Q(
        \i_iq_demod/filtre_I/tot_adder/n32 ) );
  OAI220 \i_iq_demod/filtre_I/tot_adder/U25  ( .A(
        \i_iq_demod/filtre_I/tot_adder/n31 ), .B(
        \i_iq_demod/filtre_I/tot_adder/n32 ), .C(
        \i_iq_demod/filtre_I/tot_adder/n33 ), .D(
        \i_iq_demod/filtre_I/tot_adder/n34 ), .Q(
        \i_iq_demod/filtre_I/tot_adder/n28 ) );
  NOR20 \i_iq_demod/filtre_I/tot_adder/U11  ( .A(n158), .B(n181), .Q(
        \i_iq_demod/filtre_I/tot_adder/n18 ) );
  XNR20 \i_iq_demod/filtre_I/tot_adder/U10  ( .A(
        \i_iq_demod/filtre_I/tot_adder/n17 ), .B(
        \i_iq_demod/filtre_I/tot_adder/n18 ), .Q(\i_iq_demod/filtre_I/tot [1])
         );
  XOR20 \i_iq_demod/filtre_I/tot_adder/U8  ( .A(
        \i_iq_demod/filtre_I/tot_adder/n13 ), .B(
        \i_iq_demod/filtre_I/tot_adder/n14 ), .Q(\i_iq_demod/filtre_I/tot [3])
         );
  XOR20 \i_iq_demod/filtre_I/tot_adder/U6  ( .A(
        \i_iq_demod/filtre_I/tot_adder/n9 ), .B(
        \i_iq_demod/filtre_I/tot_adder/n10 ), .Q(\i_iq_demod/filtre_I/tot [5])
         );
  XOR20 \i_iq_demod/filtre_I/tot_adder/U4  ( .A(
        \i_iq_demod/filtre_I/tot_adder/n5 ), .B(
        \i_iq_demod/filtre_I/tot_adder/n6 ), .Q(\i_iq_demod/filtre_I/tot [7])
         );
  XOR20 \i_iq_demod/filtre_I/tot_adder/U2  ( .A(
        \i_iq_demod/filtre_I/tot_adder/n1 ), .B(
        \i_iq_demod/filtre_I/tot_adder/n2 ), .Q(\i_iq_demod/filtre_I/tot [9])
         );
  NOR20 \i_iq_demod/filtre_Q/U95  ( .A(\i_iq_demod/filtre_Q/shift_count [2]), 
        .B(\i_iq_demod/filtre_Q/shift_count [0]), .Q(n1398) );
  NAND20 \i_iq_demod/filtre_Q/U40  ( .A(\i_iq_demod/filtre_Q/current_state [1]), .B(n1385), .Q(n1390) );
  OAI220 \i_iq_demod/filtre_Q/U39  ( .A(\i_iq_demod/filtre_Q/current_state [1]), .B(\i_iq_demod/filtre_Q/next_state [0]), .C(n1390), .D(
        \i_iq_demod/filtre_Q/current_state [0]), .Q(
        \i_iq_demod/filtre_Q/next_state [1]) );
  CLKIN0 \i_iq_demod/filtre_Q/U37  ( .A(n1390), .Q(n1388) );
  AOI210 \i_iq_demod/filtre_Q/U34  ( .A(\i_iq_demod/filtre_Q/current_state [2]), .B(n1387), .C(n1388), .Q(n1386) );
  DFEC1 \i_iq_demod/filtre_Q/data_out_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/temp [9]), .E(\i_iq_demod/filtre_Q/N123 ), .C(
        clk_i), .RN(resetn_i), .Q(demod_iq_qbb_o[0]) );
  DFEC1 \i_iq_demod/filtre_Q/data_out_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/temp [10]), .E(\i_iq_demod/filtre_Q/N123 ), .C(
        clk_i), .RN(resetn_i), .Q(demod_iq_qbb_o[1]) );
  DFEC1 \i_iq_demod/filtre_Q/data_out_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/temp [11]), .E(\i_iq_demod/filtre_Q/N123 ), .C(
        clk_i), .RN(resetn_i), .Q(demod_iq_qbb_o[2]) );
  DFEC1 \i_iq_demod/filtre_Q/data_out_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/temp [12]), .E(\i_iq_demod/filtre_Q/N123 ), .C(
        clk_i), .RN(resetn_i), .Q(demod_iq_qbb_o[3]) );
  DFEC1 \i_iq_demod/filtre_Q/data_out_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/temp [13]), .E(\i_iq_demod/filtre_Q/N123 ), .C(
        clk_i), .RN(resetn_i), .Q(demod_iq_qbb_o[4]) );
  DFC1 \i_iq_demod/filtre_Q/out_valid_reg  ( .D(\i_iq_demod/filtre_Q/N123 ), 
        .C(clk_i), .RN(resetn_i), .QN(n1411) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[13]  ( .D(\i_iq_demod/filtre_Q/N28 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [13]) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[12]  ( .D(\i_iq_demod/filtre_Q/N27 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [12]) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[11]  ( .D(\i_iq_demod/filtre_Q/N26 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [11]), .QN(n247)
         );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[10]  ( .D(\i_iq_demod/filtre_Q/N25 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [10]) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[9]  ( .D(\i_iq_demod/filtre_Q/N24 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [9]), .QN(n248) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[8]  ( .D(\i_iq_demod/filtre_Q/N23 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [8]) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[7]  ( .D(\i_iq_demod/filtre_Q/N22 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [7]), .QN(n239) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[6]  ( .D(\i_iq_demod/filtre_Q/N21 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [6]) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[5]  ( .D(\i_iq_demod/filtre_Q/N20 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [5]), .QN(n240) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[4]  ( .D(\i_iq_demod/filtre_Q/N19 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [4]) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[3]  ( .D(\i_iq_demod/filtre_Q/N18 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [3]), .QN(n230) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[2]  ( .D(\i_iq_demod/filtre_Q/N17 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [2]) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[1]  ( .D(\i_iq_demod/filtre_Q/N16 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/temp [1]) );
  DFC1 \i_iq_demod/filtre_Q/temp_reg[0]  ( .D(\i_iq_demod/filtre_Q/N15 ), .C(
        clk_i), .RN(resetn_i), .QN(n227) );
  DFC1 \i_iq_demod/filtre_Q/data_1_1_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/data_1_1_req [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_1_1 [4]) );
  DFC1 \i_iq_demod/filtre_Q/data_1_1_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/data_1_1_req [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_1_1 [3]) );
  DFC1 \i_iq_demod/filtre_Q/data_1_1_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/data_1_1_req [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_1_1 [2]) );
  DFC1 \i_iq_demod/filtre_Q/data_2_1_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/data_2_1_req [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_2_1 [4]) );
  DFC1 \i_iq_demod/filtre_Q/data_2_1_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/data_2_1_req [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_2_1 [3]) );
  DFC1 \i_iq_demod/filtre_Q/data_2_1_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/data_2_1_req [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_2_1 [2]) );
  DFC1 \i_iq_demod/filtre_Q/data_1_2_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/data_1_2_req [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_1_2 [4]) );
  DFC1 \i_iq_demod/filtre_Q/data_1_2_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/data_1_2_req [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_1_2 [3]) );
  DFC1 \i_iq_demod/filtre_Q/data_1_2_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/data_1_2_req [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_1_2 [2]) );
  DFC1 \i_iq_demod/filtre_Q/data_2_2_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/data_2_2_req [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_2_2 [4]) );
  DFC1 \i_iq_demod/filtre_Q/data_2_2_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/data_2_2_req [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_2_2 [3]) );
  DFC1 \i_iq_demod/filtre_Q/data_2_2_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/data_2_2_req [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_2_2 [2]), .QN(n1611) );
  DFC1 \i_iq_demod/filtre_Q/out_factor1_reg[8]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1_req [8]), .C(clk_i), .RN(resetn_i), 
        .QN(n211) );
  DFC1 \i_iq_demod/filtre_Q/out_factor1_reg[7]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1_req [7]), .C(clk_i), .RN(resetn_i), 
        .QN(n207) );
  DFC1 \i_iq_demod/filtre_Q/out_factor1_reg[6]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1_req [6]), .C(clk_i), .RN(resetn_i), 
        .QN(n155) );
  DFC1 \i_iq_demod/filtre_Q/out_factor1_reg[5]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1_req [5]), .C(clk_i), .RN(resetn_i), 
        .QN(n140) );
  DFC1 \i_iq_demod/filtre_Q/out_factor1_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1_req [0]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_Q/out_factor1 [0]), .QN(n144) );
  DFC1 \i_iq_demod/filtre_Q/out_factor2_reg[8]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2_req [4]), .C(clk_i), .RN(resetn_i), 
        .QN(n176) );
  DFC1 \i_iq_demod/filtre_Q/out_factor2_reg[7]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2_req [6]), .C(clk_i), .RN(resetn_i), 
        .QN(n172) );
  DFC1 \i_iq_demod/filtre_Q/out_factor2_reg[6]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2_req [6]), .C(clk_i), .RN(resetn_i), 
        .QN(n170) );
  DFC1 \i_iq_demod/filtre_Q/out_factor2_reg[5]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2_req [4]), .C(clk_i), .RN(resetn_i), 
        .QN(n141) );
  DFC3 \i_iq_demod/filtre_Q/current_state_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/next_state [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/current_state [1]), .QN(n1387) );
  DFC1 \i_iq_demod/filtre_Q/current_state_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/sel [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/current_state [2]), .QN(n1385) );
  DFC1 \i_iq_demod/filtre_Q/current_state_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/next_state [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/current_state [0]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U44  ( .A(
        \i_iq_demod/filtre_Q/shift_reg11 [0]), .B(n1355), .C(
        \i_iq_demod/filtre_Q/shift_reg13 [0]), .D(n1356), .Q(n1381) );
  NAND20 \i_iq_demod/filtre_Q/data_reg2/U42  ( .A(
        \i_iq_demod/filtre_Q/shift_reg15 [0]), .B(n1354), .Q(n1382) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U39  ( .A(
        \i_iq_demod/filtre_Q/shift_reg17 [0]), .B(n1352), .C(
        \i_iq_demod/filtre_Q/shift_reg19 [0]), .D(n1353), .Q(n1383) );
  NAND30 \i_iq_demod/filtre_Q/data_reg2/U38  ( .A(n1381), .B(n1382), .C(n1383), 
        .Q(\i_iq_demod/filtre_Q/data_1_2_req [0]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U37  ( .A(
        \i_iq_demod/filtre_Q/shift_reg11 [1]), .B(n1355), .C(
        \i_iq_demod/filtre_Q/shift_reg13 [1]), .D(n1356), .Q(n1378) );
  NAND20 \i_iq_demod/filtre_Q/data_reg2/U36  ( .A(
        \i_iq_demod/filtre_Q/shift_reg15 [1]), .B(n1354), .Q(n1379) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U35  ( .A(
        \i_iq_demod/filtre_Q/shift_reg17 [1]), .B(n1352), .C(
        \i_iq_demod/filtre_Q/shift_reg19 [1]), .D(n1353), .Q(n1380) );
  NAND30 \i_iq_demod/filtre_Q/data_reg2/U34  ( .A(n1378), .B(n1379), .C(n1380), 
        .Q(\i_iq_demod/filtre_Q/data_1_2_req [1]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U33  ( .A(
        \i_iq_demod/filtre_Q/shift_reg11 [2]), .B(n1355), .C(
        \i_iq_demod/filtre_Q/shift_reg13 [2]), .D(n1356), .Q(n1375) );
  NAND20 \i_iq_demod/filtre_Q/data_reg2/U32  ( .A(
        \i_iq_demod/filtre_Q/shift_reg15 [2]), .B(n1354), .Q(n1376) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U31  ( .A(
        \i_iq_demod/filtre_Q/shift_reg17 [2]), .B(n1352), .C(
        \i_iq_demod/filtre_Q/shift_reg19 [2]), .D(n1353), .Q(n1377) );
  NAND30 \i_iq_demod/filtre_Q/data_reg2/U30  ( .A(n1375), .B(n1376), .C(n1377), 
        .Q(\i_iq_demod/filtre_Q/data_1_2_req [2]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U29  ( .A(
        \i_iq_demod/filtre_Q/shift_reg11 [3]), .B(n1355), .C(
        \i_iq_demod/filtre_Q/shift_reg13 [3]), .D(n1356), .Q(n1372) );
  NAND20 \i_iq_demod/filtre_Q/data_reg2/U28  ( .A(
        \i_iq_demod/filtre_Q/shift_reg15 [3]), .B(n1354), .Q(n1373) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U27  ( .A(
        \i_iq_demod/filtre_Q/shift_reg17 [3]), .B(n1352), .C(
        \i_iq_demod/filtre_Q/shift_reg19 [3]), .D(n1353), .Q(n1374) );
  NAND30 \i_iq_demod/filtre_Q/data_reg2/U26  ( .A(n1372), .B(n1373), .C(n1374), 
        .Q(\i_iq_demod/filtre_Q/data_1_2_req [3]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U25  ( .A(
        \i_iq_demod/filtre_Q/shift_reg11 [4]), .B(n1355), .C(
        \i_iq_demod/filtre_Q/shift_reg13 [4]), .D(n1356), .Q(n1369) );
  NAND20 \i_iq_demod/filtre_Q/data_reg2/U24  ( .A(
        \i_iq_demod/filtre_Q/shift_reg15 [4]), .B(n1354), .Q(n1370) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U23  ( .A(
        \i_iq_demod/filtre_Q/shift_reg17 [4]), .B(n1352), .C(
        \i_iq_demod/filtre_Q/shift_reg19 [4]), .D(n1353), .Q(n1371) );
  NAND30 \i_iq_demod/filtre_Q/data_reg2/U22  ( .A(n1369), .B(n1370), .C(n1371), 
        .Q(\i_iq_demod/filtre_Q/data_1_2_req [4]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U21  ( .A(
        \i_iq_demod/filtre_Q/shift_reg10 [0]), .B(n1355), .C(
        \i_iq_demod/filtre_Q/shift_reg12 [0]), .D(n1356), .Q(n1366) );
  NAND20 \i_iq_demod/filtre_Q/data_reg2/U20  ( .A(
        \i_iq_demod/filtre_Q/shift_reg14 [0]), .B(n1354), .Q(n1367) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U19  ( .A(
        \i_iq_demod/filtre_Q/shift_reg16 [0]), .B(n1352), .C(
        \i_iq_demod/filtre_Q/shift_reg18 [0]), .D(n1353), .Q(n1368) );
  NAND30 \i_iq_demod/filtre_Q/data_reg2/U18  ( .A(n1366), .B(n1367), .C(n1368), 
        .Q(\i_iq_demod/filtre_Q/data_2_2_req [0]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U17  ( .A(
        \i_iq_demod/filtre_Q/shift_reg10 [1]), .B(n1355), .C(
        \i_iq_demod/filtre_Q/shift_reg12 [1]), .D(n1356), .Q(n1363) );
  NAND20 \i_iq_demod/filtre_Q/data_reg2/U16  ( .A(
        \i_iq_demod/filtre_Q/shift_reg14 [1]), .B(n1354), .Q(n1364) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U15  ( .A(
        \i_iq_demod/filtre_Q/shift_reg16 [1]), .B(n1352), .C(
        \i_iq_demod/filtre_Q/shift_reg18 [1]), .D(n1353), .Q(n1365) );
  NAND30 \i_iq_demod/filtre_Q/data_reg2/U14  ( .A(n1363), .B(n1364), .C(n1365), 
        .Q(\i_iq_demod/filtre_Q/data_2_2_req [1]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U13  ( .A(
        \i_iq_demod/filtre_Q/shift_reg10 [2]), .B(n1355), .C(
        \i_iq_demod/filtre_Q/shift_reg12 [2]), .D(n1356), .Q(n1360) );
  NAND20 \i_iq_demod/filtre_Q/data_reg2/U12  ( .A(
        \i_iq_demod/filtre_Q/shift_reg14 [2]), .B(n1354), .Q(n1361) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U11  ( .A(
        \i_iq_demod/filtre_Q/shift_reg16 [2]), .B(n1352), .C(
        \i_iq_demod/filtre_Q/shift_reg18 [2]), .D(n1353), .Q(n1362) );
  NAND30 \i_iq_demod/filtre_Q/data_reg2/U10  ( .A(n1360), .B(n1361), .C(n1362), 
        .Q(\i_iq_demod/filtre_Q/data_2_2_req [2]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U9  ( .A(
        \i_iq_demod/filtre_Q/shift_reg10 [3]), .B(n1355), .C(
        \i_iq_demod/filtre_Q/shift_reg12 [3]), .D(n1356), .Q(n1357) );
  NAND20 \i_iq_demod/filtre_Q/data_reg2/U8  ( .A(
        \i_iq_demod/filtre_Q/shift_reg14 [3]), .B(n1354), .Q(n1358) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U7  ( .A(
        \i_iq_demod/filtre_Q/shift_reg16 [3]), .B(n1352), .C(
        \i_iq_demod/filtre_Q/shift_reg18 [3]), .D(n1353), .Q(n1359) );
  NAND30 \i_iq_demod/filtre_Q/data_reg2/U6  ( .A(n1357), .B(n1358), .C(n1359), 
        .Q(\i_iq_demod/filtre_Q/data_2_2_req [3]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U5  ( .A(
        \i_iq_demod/filtre_Q/shift_reg10 [4]), .B(n1355), .C(
        \i_iq_demod/filtre_Q/shift_reg12 [4]), .D(n1356), .Q(n1349) );
  NAND20 \i_iq_demod/filtre_Q/data_reg2/U4  ( .A(
        \i_iq_demod/filtre_Q/shift_reg14 [4]), .B(n1354), .Q(n1350) );
  AOI220 \i_iq_demod/filtre_Q/data_reg2/U3  ( .A(
        \i_iq_demod/filtre_Q/shift_reg16 [4]), .B(n1352), .C(
        \i_iq_demod/filtre_Q/shift_reg18 [4]), .D(n1353), .Q(n1351) );
  NAND30 \i_iq_demod/filtre_Q/data_reg2/U2  ( .A(n1349), .B(n1350), .C(n1351), 
        .Q(\i_iq_demod/filtre_Q/data_2_2_req [4]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U44  ( .A(
        \i_iq_demod/filtre_Q/shift_reg8 [0]), .B(n1318), .C(
        \i_iq_demod/filtre_Q/shift_reg6 [0]), .D(n1319), .Q(n1344) );
  NAND20 \i_iq_demod/filtre_Q/data_reg1/U42  ( .A(
        \i_iq_demod/filtre_Q/shift_reg4 [0]), .B(n1317), .Q(n1345) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U39  ( .A(
        \i_iq_demod/filtre_Q/shift_reg2 [0]), .B(n1315), .C(
        \i_iq_demod/filtre_Q/shift_reg0 [0]), .D(n1316), .Q(n1346) );
  NAND30 \i_iq_demod/filtre_Q/data_reg1/U38  ( .A(n1344), .B(n1345), .C(n1346), 
        .Q(\i_iq_demod/filtre_Q/data_1_1_req [0]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U37  ( .A(
        \i_iq_demod/filtre_Q/shift_reg8 [1]), .B(n1318), .C(
        \i_iq_demod/filtre_Q/shift_reg6 [1]), .D(n1319), .Q(n1341) );
  NAND20 \i_iq_demod/filtre_Q/data_reg1/U36  ( .A(
        \i_iq_demod/filtre_Q/shift_reg4 [1]), .B(n1317), .Q(n1342) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U35  ( .A(
        \i_iq_demod/filtre_Q/shift_reg2 [1]), .B(n1315), .C(
        \i_iq_demod/filtre_Q/shift_reg0 [1]), .D(n1316), .Q(n1343) );
  NAND30 \i_iq_demod/filtre_Q/data_reg1/U34  ( .A(n1341), .B(n1342), .C(n1343), 
        .Q(\i_iq_demod/filtre_Q/data_1_1_req [1]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U33  ( .A(
        \i_iq_demod/filtre_Q/shift_reg8 [2]), .B(n1318), .C(
        \i_iq_demod/filtre_Q/shift_reg6 [2]), .D(n1319), .Q(n1338) );
  NAND20 \i_iq_demod/filtre_Q/data_reg1/U32  ( .A(
        \i_iq_demod/filtre_Q/shift_reg4 [2]), .B(n1317), .Q(n1339) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U31  ( .A(
        \i_iq_demod/filtre_Q/shift_reg2 [2]), .B(n1315), .C(
        \i_iq_demod/filtre_Q/shift_reg0 [2]), .D(n1316), .Q(n1340) );
  NAND30 \i_iq_demod/filtre_Q/data_reg1/U30  ( .A(n1338), .B(n1339), .C(n1340), 
        .Q(\i_iq_demod/filtre_Q/data_1_1_req [2]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U29  ( .A(
        \i_iq_demod/filtre_Q/shift_reg8 [3]), .B(n1318), .C(
        \i_iq_demod/filtre_Q/shift_reg6 [3]), .D(n1319), .Q(n1335) );
  NAND20 \i_iq_demod/filtre_Q/data_reg1/U28  ( .A(
        \i_iq_demod/filtre_Q/shift_reg4 [3]), .B(n1317), .Q(n1336) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U27  ( .A(
        \i_iq_demod/filtre_Q/shift_reg2 [3]), .B(n1315), .C(
        \i_iq_demod/filtre_Q/shift_reg0 [3]), .D(n1316), .Q(n1337) );
  NAND30 \i_iq_demod/filtre_Q/data_reg1/U26  ( .A(n1335), .B(n1336), .C(n1337), 
        .Q(\i_iq_demod/filtre_Q/data_1_1_req [3]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U25  ( .A(
        \i_iq_demod/filtre_Q/shift_reg8 [4]), .B(n1318), .C(
        \i_iq_demod/filtre_Q/shift_reg6 [4]), .D(n1319), .Q(n1332) );
  NAND20 \i_iq_demod/filtre_Q/data_reg1/U24  ( .A(
        \i_iq_demod/filtre_Q/shift_reg4 [4]), .B(n1317), .Q(n1333) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U23  ( .A(
        \i_iq_demod/filtre_Q/shift_reg2 [4]), .B(n1315), .C(
        \i_iq_demod/filtre_Q/shift_reg0 [4]), .D(n1316), .Q(n1334) );
  NAND30 \i_iq_demod/filtre_Q/data_reg1/U22  ( .A(n1332), .B(n1333), .C(n1334), 
        .Q(\i_iq_demod/filtre_Q/data_1_1_req [4]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U21  ( .A(
        \i_iq_demod/filtre_Q/shift_reg9 [0]), .B(n1318), .C(
        \i_iq_demod/filtre_Q/shift_reg7 [0]), .D(n1319), .Q(n1329) );
  NAND20 \i_iq_demod/filtre_Q/data_reg1/U20  ( .A(
        \i_iq_demod/filtre_Q/shift_reg5 [0]), .B(n1317), .Q(n1330) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U19  ( .A(
        \i_iq_demod/filtre_Q/shift_reg3 [0]), .B(n1315), .C(
        \i_iq_demod/filtre_Q/shift_reg1 [0]), .D(n1316), .Q(n1331) );
  NAND30 \i_iq_demod/filtre_Q/data_reg1/U18  ( .A(n1329), .B(n1330), .C(n1331), 
        .Q(\i_iq_demod/filtre_Q/data_2_1_req [0]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U17  ( .A(
        \i_iq_demod/filtre_Q/shift_reg9 [1]), .B(n1318), .C(
        \i_iq_demod/filtre_Q/shift_reg7 [1]), .D(n1319), .Q(n1326) );
  NAND20 \i_iq_demod/filtre_Q/data_reg1/U16  ( .A(
        \i_iq_demod/filtre_Q/shift_reg5 [1]), .B(n1317), .Q(n1327) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U15  ( .A(
        \i_iq_demod/filtre_Q/shift_reg3 [1]), .B(n1315), .C(
        \i_iq_demod/filtre_Q/shift_reg1 [1]), .D(n1316), .Q(n1328) );
  NAND30 \i_iq_demod/filtre_Q/data_reg1/U14  ( .A(n1326), .B(n1327), .C(n1328), 
        .Q(\i_iq_demod/filtre_Q/data_2_1_req [1]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U13  ( .A(
        \i_iq_demod/filtre_Q/shift_reg9 [2]), .B(n1318), .C(
        \i_iq_demod/filtre_Q/shift_reg7 [2]), .D(n1319), .Q(n1323) );
  NAND20 \i_iq_demod/filtre_Q/data_reg1/U12  ( .A(
        \i_iq_demod/filtre_Q/shift_reg5 [2]), .B(n1317), .Q(n1324) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U11  ( .A(
        \i_iq_demod/filtre_Q/shift_reg3 [2]), .B(n1315), .C(
        \i_iq_demod/filtre_Q/shift_reg1 [2]), .D(n1316), .Q(n1325) );
  NAND30 \i_iq_demod/filtre_Q/data_reg1/U10  ( .A(n1323), .B(n1324), .C(n1325), 
        .Q(\i_iq_demod/filtre_Q/data_2_1_req [2]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U9  ( .A(
        \i_iq_demod/filtre_Q/shift_reg9 [3]), .B(n1318), .C(
        \i_iq_demod/filtre_Q/shift_reg7 [3]), .D(n1319), .Q(n1320) );
  NAND20 \i_iq_demod/filtre_Q/data_reg1/U8  ( .A(
        \i_iq_demod/filtre_Q/shift_reg5 [3]), .B(n1317), .Q(n1321) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U7  ( .A(
        \i_iq_demod/filtre_Q/shift_reg3 [3]), .B(n1315), .C(
        \i_iq_demod/filtre_Q/shift_reg1 [3]), .D(n1316), .Q(n1322) );
  NAND30 \i_iq_demod/filtre_Q/data_reg1/U6  ( .A(n1320), .B(n1321), .C(n1322), 
        .Q(\i_iq_demod/filtre_Q/data_2_1_req [3]) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U5  ( .A(
        \i_iq_demod/filtre_Q/shift_reg9 [4]), .B(n1318), .C(
        \i_iq_demod/filtre_Q/shift_reg7 [4]), .D(n1319), .Q(n1312) );
  NAND20 \i_iq_demod/filtre_Q/data_reg1/U4  ( .A(
        \i_iq_demod/filtre_Q/shift_reg5 [4]), .B(n1317), .Q(n1313) );
  AOI220 \i_iq_demod/filtre_Q/data_reg1/U3  ( .A(
        \i_iq_demod/filtre_Q/shift_reg3 [4]), .B(n1315), .C(
        \i_iq_demod/filtre_Q/shift_reg1 [4]), .D(n1316), .Q(n1314) );
  NAND30 \i_iq_demod/filtre_Q/data_reg1/U2  ( .A(n1312), .B(n1313), .C(n1314), 
        .Q(\i_iq_demod/filtre_Q/data_2_1_req [4]) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U44  ( .A(
        \i_iq_demod/filtre_I/shift_reg11 [0]), .B(n1282), .C(
        \i_iq_demod/filtre_I/shift_reg13 [0]), .D(n1283), .Q(n1308) );
  NAND20 \i_iq_demod/filtre_I/data_reg2/U42  ( .A(
        \i_iq_demod/filtre_I/shift_reg15 [0]), .B(n1281), .Q(n1309) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U39  ( .A(
        \i_iq_demod/filtre_I/shift_reg17 [0]), .B(n1279), .C(
        \i_iq_demod/filtre_I/shift_reg19 [0]), .D(n1280), .Q(n1310) );
  NAND30 \i_iq_demod/filtre_I/data_reg2/U38  ( .A(n1308), .B(n1309), .C(n1310), 
        .Q(\i_iq_demod/filtre_I/data_1_2_req [0]) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U37  ( .A(
        \i_iq_demod/filtre_I/shift_reg11 [1]), .B(n1282), .C(
        \i_iq_demod/filtre_I/shift_reg13 [1]), .D(n1283), .Q(n1305) );
  NAND20 \i_iq_demod/filtre_I/data_reg2/U36  ( .A(
        \i_iq_demod/filtre_I/shift_reg15 [1]), .B(n1281), .Q(n1306) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U35  ( .A(
        \i_iq_demod/filtre_I/shift_reg17 [1]), .B(n1279), .C(
        \i_iq_demod/filtre_I/shift_reg19 [1]), .D(n1280), .Q(n1307) );
  NAND30 \i_iq_demod/filtre_I/data_reg2/U34  ( .A(n1305), .B(n1306), .C(n1307), 
        .Q(\i_iq_demod/filtre_I/data_1_2_req [1]) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U33  ( .A(
        \i_iq_demod/filtre_I/shift_reg11 [2]), .B(n1282), .C(
        \i_iq_demod/filtre_I/shift_reg13 [2]), .D(n1283), .Q(n1302) );
  NAND20 \i_iq_demod/filtre_I/data_reg2/U32  ( .A(
        \i_iq_demod/filtre_I/shift_reg15 [2]), .B(n1281), .Q(n1303) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U31  ( .A(
        \i_iq_demod/filtre_I/shift_reg17 [2]), .B(n1279), .C(
        \i_iq_demod/filtre_I/shift_reg19 [2]), .D(n1280), .Q(n1304) );
  NAND30 \i_iq_demod/filtre_I/data_reg2/U30  ( .A(n1302), .B(n1303), .C(n1304), 
        .Q(\i_iq_demod/filtre_I/data_1_2_req [2]) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U29  ( .A(
        \i_iq_demod/filtre_I/shift_reg11 [3]), .B(n1282), .C(
        \i_iq_demod/filtre_I/shift_reg13 [3]), .D(n1283), .Q(n1299) );
  NAND20 \i_iq_demod/filtre_I/data_reg2/U28  ( .A(
        \i_iq_demod/filtre_I/shift_reg15 [3]), .B(n1281), .Q(n1300) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U27  ( .A(
        \i_iq_demod/filtre_I/shift_reg17 [3]), .B(n1279), .C(
        \i_iq_demod/filtre_I/shift_reg19 [3]), .D(n1280), .Q(n1301) );
  NAND30 \i_iq_demod/filtre_I/data_reg2/U26  ( .A(n1299), .B(n1300), .C(n1301), 
        .Q(\i_iq_demod/filtre_I/data_1_2_req [3]) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U25  ( .A(
        \i_iq_demod/filtre_I/shift_reg11 [4]), .B(n1282), .C(
        \i_iq_demod/filtre_I/shift_reg13 [4]), .D(n1283), .Q(n1296) );
  NAND20 \i_iq_demod/filtre_I/data_reg2/U24  ( .A(
        \i_iq_demod/filtre_I/shift_reg15 [4]), .B(n1281), .Q(n1297) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U23  ( .A(
        \i_iq_demod/filtre_I/shift_reg17 [4]), .B(n1279), .C(
        \i_iq_demod/filtre_I/shift_reg19 [4]), .D(n1280), .Q(n1298) );
  NAND30 \i_iq_demod/filtre_I/data_reg2/U22  ( .A(n1296), .B(n1297), .C(n1298), 
        .Q(\i_iq_demod/filtre_I/data_1_2_req [4]) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U21  ( .A(
        \i_iq_demod/filtre_I/shift_reg10 [0]), .B(n1282), .C(
        \i_iq_demod/filtre_I/shift_reg12 [0]), .D(n1283), .Q(n1293) );
  NAND20 \i_iq_demod/filtre_I/data_reg2/U20  ( .A(
        \i_iq_demod/filtre_I/shift_reg14 [0]), .B(n1281), .Q(n1294) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U19  ( .A(
        \i_iq_demod/filtre_I/shift_reg16 [0]), .B(n1279), .C(
        \i_iq_demod/filtre_I/shift_reg18 [0]), .D(n1280), .Q(n1295) );
  NAND30 \i_iq_demod/filtre_I/data_reg2/U18  ( .A(n1293), .B(n1294), .C(n1295), 
        .Q(\i_iq_demod/filtre_I/data_2_2_req [0]) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U17  ( .A(
        \i_iq_demod/filtre_I/shift_reg10 [1]), .B(n1282), .C(
        \i_iq_demod/filtre_I/shift_reg12 [1]), .D(n1283), .Q(n1290) );
  NAND20 \i_iq_demod/filtre_I/data_reg2/U16  ( .A(
        \i_iq_demod/filtre_I/shift_reg14 [1]), .B(n1281), .Q(n1291) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U15  ( .A(
        \i_iq_demod/filtre_I/shift_reg16 [1]), .B(n1279), .C(
        \i_iq_demod/filtre_I/shift_reg18 [1]), .D(n1280), .Q(n1292) );
  NAND30 \i_iq_demod/filtre_I/data_reg2/U14  ( .A(n1290), .B(n1291), .C(n1292), 
        .Q(\i_iq_demod/filtre_I/data_2_2_req [1]) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U13  ( .A(
        \i_iq_demod/filtre_I/shift_reg10 [2]), .B(n1282), .C(
        \i_iq_demod/filtre_I/shift_reg12 [2]), .D(n1283), .Q(n1287) );
  NAND20 \i_iq_demod/filtre_I/data_reg2/U12  ( .A(
        \i_iq_demod/filtre_I/shift_reg14 [2]), .B(n1281), .Q(n1288) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U11  ( .A(
        \i_iq_demod/filtre_I/shift_reg16 [2]), .B(n1279), .C(
        \i_iq_demod/filtre_I/shift_reg18 [2]), .D(n1280), .Q(n1289) );
  NAND30 \i_iq_demod/filtre_I/data_reg2/U10  ( .A(n1287), .B(n1288), .C(n1289), 
        .Q(\i_iq_demod/filtre_I/data_2_2_req [2]) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U9  ( .A(
        \i_iq_demod/filtre_I/shift_reg10 [3]), .B(n1282), .C(
        \i_iq_demod/filtre_I/shift_reg12 [3]), .D(n1283), .Q(n1284) );
  NAND20 \i_iq_demod/filtre_I/data_reg2/U8  ( .A(
        \i_iq_demod/filtre_I/shift_reg14 [3]), .B(n1281), .Q(n1285) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U7  ( .A(
        \i_iq_demod/filtre_I/shift_reg16 [3]), .B(n1279), .C(
        \i_iq_demod/filtre_I/shift_reg18 [3]), .D(n1280), .Q(n1286) );
  NAND30 \i_iq_demod/filtre_I/data_reg2/U6  ( .A(n1284), .B(n1285), .C(n1286), 
        .Q(\i_iq_demod/filtre_I/data_2_2_req [3]) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U5  ( .A(
        \i_iq_demod/filtre_I/shift_reg10 [4]), .B(n1282), .C(
        \i_iq_demod/filtre_I/shift_reg12 [4]), .D(n1283), .Q(n1276) );
  NAND20 \i_iq_demod/filtre_I/data_reg2/U4  ( .A(
        \i_iq_demod/filtre_I/shift_reg14 [4]), .B(n1281), .Q(n1277) );
  AOI220 \i_iq_demod/filtre_I/data_reg2/U3  ( .A(
        \i_iq_demod/filtre_I/shift_reg16 [4]), .B(n1279), .C(
        \i_iq_demod/filtre_I/shift_reg18 [4]), .D(n1280), .Q(n1278) );
  NAND30 \i_iq_demod/filtre_I/data_reg2/U2  ( .A(n1276), .B(n1277), .C(n1278), 
        .Q(\i_iq_demod/filtre_I/data_2_2_req [4]) );
  NOR30 \i_iq_demod/filtre_Q/factor/U80  ( .A(\i_iq_demod/filtre_Q/sel [0]), 
        .B(\i_iq_demod/filtre_Q/sel [1]), .C(n1348), .Q(n1266) );
  NOR30 \i_iq_demod/filtre_Q/factor/U75  ( .A(\i_iq_demod/filtre_Q/sel [0]), 
        .B(n1944), .C(n1389), .Q(n1265) );
  NAND20 \i_iq_demod/filtre_Q/shift_r/U9  ( .A(
        \i_iq_demod/filtre_Q/shift_count [0]), .B(
        \i_iq_demod/filtre_Q/shift_count [1]), .Q(n1261) );
  XNR20 \i_iq_demod/filtre_Q/shift_r/U7  ( .A(n1258), .B(
        \i_iq_demod/filtre_Q/shift_count [0]), .Q(
        \i_iq_demod/filtre_Q/shift_r/N9 ) );
  AOI210 \i_iq_demod/filtre_Q/shift_r/U6  ( .A(n1261), .B(
        \i_iq_demod/demod/validation/n3 ), .C(\i_iq_demod/filtre_Q/shift_r/N9 ), .Q(n1262) );
  CLKIN0 \i_iq_demod/filtre_Q/shift_r/U5  ( .A(n1261), .Q(n1259) );
  NOR40 \i_iq_demod/filtre_Q/shift_r/U4  ( .A(n1259), .B(
        \i_iq_demod/filtre_Q/shift_r/N9 ), .C(n1260), .D(
        \i_iq_demod/demod/validation/n3 ), .Q(\i_iq_demod/filtre_Q/shift_r/N3 ) );
  AOI310 \i_iq_demod/filtre_Q/shift_r/U3  ( .A(
        \i_iq_demod/filtre_Q/shift_count [2]), .B(n1258), .C(
        \i_iq_demod/filter_en ), .D(\i_iq_demod/filtre_Q/shift_count [0]), .Q(
        \i_iq_demod/filtre_Q/shift_r/N8 ) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out19_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg18 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg19 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out18_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg17 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg18 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out17_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg16 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg17 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out16_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg15 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg16 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out15_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg14 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg15 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out14_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg13 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg14 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out13_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg12 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg13 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out12_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg11 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg12 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out11_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg10 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg11 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out10_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg9 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg10 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out9_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg8 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg9 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out8_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg7 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg8 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out7_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg6 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg7 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out6_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg5 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg6 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out5_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg4 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg5 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out4_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg3 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg4 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out3_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg2 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg3 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out2_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg1 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg2 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out1_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg0 [0]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg1 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out0_reg[0]  ( .D(
        \i_iq_demod/Q_BB_IN [0]), .E(n266), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/shift_reg0 [0]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out19_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg18 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg19 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out18_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg17 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg18 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out17_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg16 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg17 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out16_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg15 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg16 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out15_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg14 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg15 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out14_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg13 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg14 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out13_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg12 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg13 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out12_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg11 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg12 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out11_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg10 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg11 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out10_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg9 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg10 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out9_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg8 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg9 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out8_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg7 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg8 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out7_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg6 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg7 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out6_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg5 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg6 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out5_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg4 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg5 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out4_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg3 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg4 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out3_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg2 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg3 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out2_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg1 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg2 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out1_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg0 [1]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg1 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out0_reg[1]  ( .D(
        \i_iq_demod/Q_BB_IN [1]), .E(n266), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/shift_reg0 [1]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out19_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg18 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg19 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out18_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg17 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg18 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out17_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg16 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg17 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out16_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg15 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg16 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out15_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg14 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg15 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out14_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg13 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg14 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out13_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg12 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg13 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out12_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg11 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg12 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out11_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg10 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg11 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out10_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg9 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg10 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out9_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg8 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg9 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out8_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg7 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg8 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out7_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg6 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg7 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out6_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg5 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg6 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out5_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg4 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg5 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out4_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg3 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg4 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out3_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg2 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg3 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out2_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg1 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg2 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out1_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg0 [2]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg1 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out0_reg[2]  ( .D(
        \i_iq_demod/Q_BB_IN [2]), .E(n266), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/shift_reg0 [2]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out19_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg18 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg19 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out18_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg17 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg18 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out17_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg16 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg17 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out16_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg15 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg16 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out15_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg14 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg15 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out14_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg13 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg14 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out13_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg12 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg13 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out12_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg11 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg12 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out11_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg10 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg11 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out10_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg9 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg10 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out9_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg8 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg9 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out8_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg7 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg8 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out7_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg6 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg7 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out6_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg5 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg6 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out5_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg4 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg5 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out4_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg3 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg4 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out3_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg2 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg3 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out2_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg1 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg2 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out1_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg0 [3]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg1 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out0_reg[3]  ( .D(
        \i_iq_demod/Q_BB_IN [3]), .E(n266), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/shift_reg0 [3]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out19_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg18 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg19 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out18_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg17 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg18 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out17_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg16 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg17 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out16_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg15 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg16 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out15_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg14 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg15 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out14_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg13 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg14 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out13_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg12 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg13 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out12_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg11 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg12 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out11_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg10 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg11 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out10_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg9 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg10 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out9_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg8 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg9 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out8_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg7 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg8 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out7_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg6 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg7 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out6_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg5 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg6 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out5_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg4 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg5 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out4_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg3 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg4 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out3_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg2 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg3 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out2_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg1 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg2 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out1_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/shift_reg0 [4]), .E(n266), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/shift_reg1 [4]) );
  DFEC1 \i_iq_demod/filtre_Q/shift_r/data_out0_reg[4]  ( .D(
        \i_iq_demod/Q_BB_IN [4]), .E(n266), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/shift_reg0 [4]) );
  JKC1 \i_iq_demod/filtre_Q/shift_r/cpt_shift_reg[2]  ( .J(n1259), .K(n1262), 
        .C(clk_i), .RN(resetn_i), .Q(\i_iq_demod/filtre_Q/shift_count [2]), 
        .QN(n1260) );
  TFEC3 \i_iq_demod/filtre_Q/shift_r/cpt_shift_reg[1]  ( .T(
        \i_iq_demod/filtre_Q/shift_count [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/shift_count [1]), .QN(n1258) );
  DFC1 \i_iq_demod/filtre_Q/shift_r/cpt_shift_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/shift_r/N8 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/shift_count [0]) );
  XNR20 \i_iq_demod/filtre_Q/temp_adder/U75  ( .A(n227), .B(
        \i_iq_demod/filtre_Q/tot [0]), .Q(\i_iq_demod/filtre_Q/n_temp [0]) );
  CLKIN0 \i_iq_demod/filtre_Q/temp_adder/U74  ( .A(
        \i_iq_demod/filtre_Q/tot [9]), .Q(n1253) );
  CLKIN0 \i_iq_demod/filtre_Q/temp_adder/U72  ( .A(
        \i_iq_demod/filtre_Q/tot [7]), .Q(n1254) );
  CLKIN0 \i_iq_demod/filtre_Q/temp_adder/U70  ( .A(
        \i_iq_demod/filtre_Q/tot [5]), .Q(n1255) );
  CLKIN0 \i_iq_demod/filtre_Q/temp_adder/U68  ( .A(
        \i_iq_demod/filtre_Q/tot [3]), .Q(n1256) );
  CLKIN0 \i_iq_demod/filtre_Q/temp_adder/U66  ( .A(
        \i_iq_demod/filtre_Q/tot [0]), .Q(n1244) );
  XNR20 \i_iq_demod/filtre_Q/temp_adder/U65  ( .A(\i_iq_demod/filtre_Q/tot [1]), .B(\i_iq_demod/filtre_Q/temp [1]), .Q(n1242) );
  NAND20 \i_iq_demod/filtre_Q/temp_adder/U64  ( .A(
        \i_iq_demod/filtre_Q/temp [1]), .B(\i_iq_demod/filtre_Q/tot [1]), .Q(
        n1257) );
  OAI310 \i_iq_demod/filtre_Q/temp_adder/U63  ( .A(n1244), .B(n1242), .C(n227), 
        .D(n1257), .Q(n1240) );
  XNR20 \i_iq_demod/filtre_Q/temp_adder/U59  ( .A(\i_iq_demod/filtre_Q/tot [3]), .B(\i_iq_demod/filtre_Q/temp [3]), .Q(n1239) );
  OAI220 \i_iq_demod/filtre_Q/temp_adder/U58  ( .A(n1256), .B(n230), .C(n1238), 
        .D(n1239), .Q(n1236) );
  XNR20 \i_iq_demod/filtre_Q/temp_adder/U54  ( .A(\i_iq_demod/filtre_Q/tot [5]), .B(\i_iq_demod/filtre_Q/temp [5]), .Q(n1235) );
  OAI220 \i_iq_demod/filtre_Q/temp_adder/U53  ( .A(n1255), .B(n240), .C(n1234), 
        .D(n1235), .Q(n1232) );
  XNR20 \i_iq_demod/filtre_Q/temp_adder/U49  ( .A(\i_iq_demod/filtre_Q/tot [7]), .B(\i_iq_demod/filtre_Q/temp [7]), .Q(n1231) );
  OAI220 \i_iq_demod/filtre_Q/temp_adder/U48  ( .A(n1254), .B(n239), .C(n1230), 
        .D(n1231), .Q(n1228) );
  XNR20 \i_iq_demod/filtre_Q/temp_adder/U44  ( .A(\i_iq_demod/filtre_Q/tot [9]), .B(\i_iq_demod/filtre_Q/temp [9]), .Q(n1227) );
  OAI220 \i_iq_demod/filtre_Q/temp_adder/U43  ( .A(n1253), .B(n248), .C(n1226), 
        .D(n1227), .Q(n1251) );
  XNR20 \i_iq_demod/filtre_Q/temp_adder/U38  ( .A(
        \i_iq_demod/filtre_Q/tot [11]), .B(\i_iq_demod/filtre_Q/temp [11]), 
        .Q(n1250) );
  XOR20 \i_iq_demod/filtre_Q/temp_adder/U37  ( .A(n1249), .B(n1250), .Q(
        \i_iq_demod/filtre_Q/n_temp [11]) );
  CLKIN0 \i_iq_demod/filtre_Q/temp_adder/U36  ( .A(
        \i_iq_demod/filtre_Q/tot [11]), .Q(n1248) );
  OAI220 \i_iq_demod/filtre_Q/temp_adder/U34  ( .A(n1248), .B(n247), .C(n1249), 
        .D(n1250), .Q(n1246) );
  NOR20 \i_iq_demod/filtre_Q/temp_adder/U11  ( .A(n227), .B(n1244), .Q(n1243)
         );
  XNR20 \i_iq_demod/filtre_Q/temp_adder/U10  ( .A(n1242), .B(n1243), .Q(
        \i_iq_demod/filtre_Q/n_temp [1]) );
  XOR20 \i_iq_demod/filtre_Q/temp_adder/U8  ( .A(n1238), .B(n1239), .Q(
        \i_iq_demod/filtre_Q/n_temp [3]) );
  XOR20 \i_iq_demod/filtre_Q/temp_adder/U6  ( .A(n1234), .B(n1235), .Q(
        \i_iq_demod/filtre_Q/n_temp [5]) );
  XOR20 \i_iq_demod/filtre_Q/temp_adder/U4  ( .A(n1230), .B(n1231), .Q(
        \i_iq_demod/filtre_Q/n_temp [7]) );
  XOR20 \i_iq_demod/filtre_Q/temp_adder/U2  ( .A(n1226), .B(n1227), .Q(
        \i_iq_demod/filtre_Q/n_temp [9]) );
  XOR20 \i_iq_demod/filtre_Q/sum2_adder/U10  ( .A(
        \i_iq_demod/filtre_Q/data_2_2 [3]), .B(
        \i_iq_demod/filtre_Q/data_1_2 [3]), .Q(n1219) );
  CLKIN0 \i_iq_demod/filtre_Q/sum2_adder/U8  ( .A(n1220), .Q(n1218) );
  XOR20 \i_iq_demod/filtre_Q/sum1_adder/U10  ( .A(
        \i_iq_demod/filtre_Q/data_2_1 [3]), .B(
        \i_iq_demod/filtre_Q/data_1_1 [3]), .Q(n1210) );
  AOI220 \i_iq_demod/filtre_Q/sum1_adder/U7  ( .A(
        \i_iq_demod/filtre_Q/data_2_1 [3]), .B(
        \i_iq_demod/filtre_Q/data_1_1 [3]), .C(n1209), .D(n1210), .Q(n1208) );
  XOR20 \i_iq_demod/filtre_I/sum2_adder/U10  ( .A(
        \i_iq_demod/filtre_I/data_2_2 [3]), .B(
        \i_iq_demod/filtre_I/data_1_2 [3]), .Q(n1201) );
  AOI220 \i_iq_demod/filtre_I/sum2_adder/U7  ( .A(
        \i_iq_demod/filtre_I/data_2_2 [3]), .B(
        \i_iq_demod/filtre_I/data_1_2 [3]), .C(n1200), .D(n1201), .Q(n1199) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U117  ( .A(n145), .B(n1770), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[0] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U107  ( .A(n141), .B(n1771), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[5] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U105  ( .A(n170), .B(n1770), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U103  ( .A(n172), .B(n1771), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[1][6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U101  ( .A(n1770), .B(n176), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[1][7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U99  ( .A(n145), .B(n210), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[0] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U96  ( .A(n128), .B(n210), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[3] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U94  ( .A(n141), .B(n210), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[5] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U92  ( .A(n172), .B(n210), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U91  ( .A(n210), .B(n176), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[9] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U88  ( .A(n153), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[1] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U85  ( .A(n151), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[4] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U84  ( .A(n141), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[5] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U83  ( .A(n170), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U82  ( .A(n172), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U81  ( .A(n1198), .B(n176), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[9] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U77  ( .A(n152), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[2] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U75  ( .A(n151), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[4] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U73  ( .A(n170), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U72  ( .A(n172), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U68  ( .A(n153), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[1] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U67  ( .A(n152), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[2] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U66  ( .A(n128), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[3] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U65  ( .A(n151), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[4] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U63  ( .A(n170), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U57  ( .A(n152), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[2] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U55  ( .A(n151), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[4] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U54  ( .A(n141), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[5] ) );
  NAND20 \i_iq_demod/filtre_Q/mult2_multiplier/U46  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe [2]), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/B_pipe ), .Q(n1196) );
  CLKIN0 \i_iq_demod/filtre_Q/mult2_multiplier/U45  ( .A(n1196), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[2] ) );
  NAND20 \i_iq_demod/filtre_Q/mult2_multiplier/U44  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe [3]), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/B_pipe ), .Q(n1195) );
  CLKIN0 \i_iq_demod/filtre_Q/mult2_multiplier/U43  ( .A(n1195), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[3] ) );
  NAND20 \i_iq_demod/filtre_Q/mult2_multiplier/U42  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe [4]), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/B_pipe ), .Q(n1194) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U24  ( .A(n172), .B(n1766), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U14  ( .A(n172), .B(n1671), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U13  ( .A(n1671), .B(n176), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[9] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U11  ( .A(n206), .B(n145), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[0] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U9  ( .A(n206), .B(n152), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[2] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U8  ( .A(n206), .B(n128), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[3] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U7  ( .A(n206), .B(n151), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[4] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U6  ( .A(n206), .B(n141), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[5] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U5  ( .A(n206), .B(n170), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U4  ( .A(n206), .B(n172), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/U3  ( .A(n206), .B(n176), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[9] ) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/B_pipe_reg  ( .D(
        \i_iq_demod/filtre_Q/_16_net_[8] ), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/B_pipe ), .QN(n96) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2 [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe [0]) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2 [1]), .C(clk_i), .RN(resetn_i), .QN(
        n95) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2 [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe [2]) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2 [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe [3]) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2 [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/A_pipe [4]) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe_reg[9][0]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[9][0] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][0] ), .QN(n217)
         );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe_reg[9][1]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[9][1] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][1] ) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe_reg[9][2]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[9][2] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][2] ) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe_reg[9][3]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[9][3] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][3] ), .QN(n222)
         );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe_reg[9][4]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[9][4] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][4] ) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/S_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[0] ), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult2 [0]), .QN(n180) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/S_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [1]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult2 [1]) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/S_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [2]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult2 [2]) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/S_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [3]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult2 [3]), .QN(n223) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/S_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [4]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult2 [4]) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/S_reg[5]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [5]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult2 [5]), .QN(n233) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/S_reg[6]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [6]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult2 [6]) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/S_reg[7]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [7]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult2 [7]), .QN(n232) );
  DFC1 \i_iq_demod/filtre_Q/mult2_multiplier/S_reg[8]  ( .D(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [8]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult2 [8]) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U117  ( .A(n144), .B(n1729), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[0] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U107  ( .A(n140), .B(n1729), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[5] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U105  ( .A(n155), .B(n1728), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U103  ( .A(n207), .B(n1728), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[1][6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U101  ( .A(n136), .B(n211), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[1][7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U97  ( .A(n199), .B(n173), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[2] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U96  ( .A(n127), .B(n173), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[3] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U95  ( .A(n150), .B(n173), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[4] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U94  ( .A(n140), .B(n173), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[5] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U93  ( .A(n155), .B(n173), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U92  ( .A(n207), .B(n173), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U91  ( .A(n173), .B(n211), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[9] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U89  ( .A(n144), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[0] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U88  ( .A(n200), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[1] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U86  ( .A(n127), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[3] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U85  ( .A(n150), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[4] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U84  ( .A(n140), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[5] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U83  ( .A(n155), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U82  ( .A(n207), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U81  ( .A(n1193), .B(n211), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[9] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U77  ( .A(n199), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[2] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U72  ( .A(n207), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U57  ( .A(n199), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[2] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U56  ( .A(n127), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[3] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U55  ( .A(n150), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[4] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U54  ( .A(n140), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[5] ) );
  NAND20 \i_iq_demod/filtre_Q/mult1_multiplier/U48  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe [1]), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/B_pipe ), .Q(n1191) );
  NAND20 \i_iq_demod/filtre_Q/mult1_multiplier/U46  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe [2]), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/B_pipe ), .Q(n1190) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/U45  ( .A(n1190), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[2] ) );
  NAND20 \i_iq_demod/filtre_Q/mult1_multiplier/U44  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe [3]), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/B_pipe ), .Q(n1189) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/U43  ( .A(n1189), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[3] ) );
  NAND20 \i_iq_demod/filtre_Q/mult1_multiplier/U42  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe [4]), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/B_pipe ), .Q(n1188) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U17  ( .A(n150), .B(n1890), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[4] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U16  ( .A(n140), .B(n1890), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[5] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U15  ( .A(n155), .B(n1890), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U14  ( .A(n207), .B(n1890), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U13  ( .A(n1890), .B(n211), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[9] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U11  ( .A(n167), .B(n144), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[0] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U10  ( .A(n167), .B(n200), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[1] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U9  ( .A(n167), .B(n199), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[2] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U8  ( .A(n167), .B(n127), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[3] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U7  ( .A(n1635), .B(n150), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[4] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U6  ( .A(n1635), .B(n140), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[5] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U5  ( .A(n1635), .B(n155), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[6] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U4  ( .A(n1635), .B(n207), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[7] ) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/U3  ( .A(n1635), .B(n211), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[9] ) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/B_pipe_reg  ( .D(
        \i_iq_demod/filtre_Q/_15_net_[8] ), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/B_pipe ) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1 [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe [0]) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1 [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe [1]) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1 [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe [2]) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1 [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe [3]) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1 [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/A_pipe [4]) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe_reg[9][0]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[9][0] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][0] ), .QN(n216)
         );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe_reg[9][1]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[9][1] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][1] ) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe_reg[9][2]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[9][2] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][2] ) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe_reg[9][3]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[9][3] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][3] ), .QN(n221)
         );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe_reg[9][4]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[9][4] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][4] ) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/S_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[0] ), .C(clk_i), .RN(
        resetn_i), .QN(n157) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/S_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [1]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult1 [1]) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/S_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [2]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult1 [2]) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/S_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [3]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult1 [3]), .QN(n183) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/S_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [4]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult1 [4]) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/S_reg[5]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [5]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult1 [5]), .QN(n188) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/S_reg[6]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [6]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult1 [6]) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/S_reg[7]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [7]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult1 [7]), .QN(n187) );
  DFC1 \i_iq_demod/filtre_Q/mult1_multiplier/S_reg[8]  ( .D(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [8]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_Q/mult1 [8]) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U107  ( .A(n139), .B(n135), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[5] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U105  ( .A(n169), .B(n135), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[6] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U103  ( .A(n171), .B(n135), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[1][6] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U101  ( .A(n135), .B(n175), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[1][7] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U98  ( .A(n149), .B(n209), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[1] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U96  ( .A(n131), .B(n209), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[3] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U95  ( .A(n147), .B(n209), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[4] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U94  ( .A(n139), .B(n209), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[5] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U93  ( .A(n169), .B(n209), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[6] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U92  ( .A(n171), .B(n209), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[7] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U91  ( .A(n209), .B(n175), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[9] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U88  ( .A(n149), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[1] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U87  ( .A(n148), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[2] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U86  ( .A(n131), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[3] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U84  ( .A(n139), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[5] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U83  ( .A(n169), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[6] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U82  ( .A(n171), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[7] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U81  ( .A(n1187), .B(n175), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[9] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U77  ( .A(n148), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[2] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U73  ( .A(n169), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[6] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U72  ( .A(n171), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[7] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U68  ( .A(n149), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[1] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U67  ( .A(n148), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[2] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U63  ( .A(n169), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[6] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U57  ( .A(n148), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[2] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U56  ( .A(n131), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[3] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U55  ( .A(n147), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[4] ) );
  NAND20 \i_iq_demod/filtre_I/mult2_multiplier/U46  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/A_pipe [2]), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/B_pipe ), .Q(n1185) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/U45  ( .A(n1185), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[2] ) );
  NAND20 \i_iq_demod/filtre_I/mult2_multiplier/U44  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/A_pipe [3]), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/B_pipe ), .Q(n1184) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/U43  ( .A(n1184), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[3] ) );
  NAND20 \i_iq_demod/filtre_I/mult2_multiplier/U42  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/A_pipe [4]), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/B_pipe ), .Q(n1183) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U27  ( .A(n147), .B(n193), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[4] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U26  ( .A(n139), .B(n193), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[5] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U24  ( .A(n171), .B(n193), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[7] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U23  ( .A(n193), .B(n175), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[9] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U17  ( .A(n147), .B(n203), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[4] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U16  ( .A(n139), .B(n203), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[5] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U15  ( .A(n169), .B(n203), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[6] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U14  ( .A(n171), .B(n203), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[7] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U13  ( .A(n203), .B(n175), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[9] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U11  ( .A(n205), .B(n143), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[0] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U8  ( .A(n205), .B(n131), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[3] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U7  ( .A(n205), .B(n147), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[4] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U6  ( .A(n205), .B(n139), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[5] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U5  ( .A(n205), .B(n169), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[6] ) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/U4  ( .A(n205), .B(n171), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[7] ) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/B_pipe_reg  ( .D(
        \i_iq_demod/filtre_I/_16_net_[8] ), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/B_pipe ), .QN(n98) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/A_pipe_reg[0]  ( .D(
        \i_iq_demod/filtre_I/out_factor2 [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/A_pipe [0]) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/A_pipe_reg[1]  ( .D(
        \i_iq_demod/filtre_I/out_factor2 [1]), .C(clk_i), .RN(resetn_i), .QN(
        n97) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/A_pipe_reg[2]  ( .D(
        \i_iq_demod/filtre_I/out_factor2 [2]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/A_pipe [2]) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/A_pipe_reg[3]  ( .D(
        \i_iq_demod/filtre_I/out_factor2 [3]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/A_pipe [3]) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/A_pipe_reg[4]  ( .D(
        \i_iq_demod/filtre_I/out_factor2 [4]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/A_pipe [4]) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/register_pipe_reg[9][0]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/register[9][0] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][0] ), .QN(n215)
         );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/register_pipe_reg[9][1]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/register[9][1] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][1] ) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/register_pipe_reg[9][2]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/register[9][2] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][2] ) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/register_pipe_reg[9][3]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/register[9][3] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][3] ), .QN(n220)
         );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/register_pipe_reg[9][4]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/register[9][4] ), .C(clk_i), 
        .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][4] ) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/S_reg[0]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[0] ), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult2 [0]), .QN(n181) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/S_reg[1]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [1]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult2 [1]) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/S_reg[2]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [2]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult2 [2]) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/S_reg[3]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [3]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult2 [3]), .QN(n224) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/S_reg[4]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [4]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult2 [4]) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/S_reg[5]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [5]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult2 [5]), .QN(n235) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/S_reg[6]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [6]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult2 [6]) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/S_reg[7]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [7]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult2 [7]), .QN(n234) );
  DFC1 \i_iq_demod/filtre_I/mult2_multiplier/S_reg[8]  ( .D(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [8]), .C(clk_i), .RN(
        resetn_i), .Q(\i_iq_demod/filtre_I/mult2 [8]) );
  XNR20 \i_iq_demod/filtre_Q/tot_adder/U66  ( .A(n157), .B(
        \i_iq_demod/filtre_Q/mult2 [0]), .Q(\i_iq_demod/filtre_Q/tot [0]) );
  CLKIN0 \i_iq_demod/filtre_Q/tot_adder/U65  ( .A(
        \i_iq_demod/filtre_Q/mult2 [9]), .Q(n1180) );
  CLKIN0 \i_iq_demod/filtre_Q/tot_adder/U64  ( .A(
        \i_iq_demod/filtre_Q/mult1 [9]), .Q(n1181) );
  XNR20 \i_iq_demod/filtre_Q/tot_adder/U56  ( .A(
        \i_iq_demod/filtre_Q/mult2 [1]), .B(\i_iq_demod/filtre_Q/mult1 [1]), 
        .Q(n1168) );
  NAND20 \i_iq_demod/filtre_Q/tot_adder/U55  ( .A(
        \i_iq_demod/filtre_Q/mult1 [1]), .B(\i_iq_demod/filtre_Q/mult2 [1]), 
        .Q(n1182) );
  OAI310 \i_iq_demod/filtre_Q/tot_adder/U54  ( .A(n180), .B(n1168), .C(n157), 
        .D(n1182), .Q(n1166) );
  XNR20 \i_iq_demod/filtre_Q/tot_adder/U50  ( .A(
        \i_iq_demod/filtre_Q/mult2 [3]), .B(\i_iq_demod/filtre_Q/mult1 [3]), 
        .Q(n1165) );
  OAI220 \i_iq_demod/filtre_Q/tot_adder/U49  ( .A(n223), .B(n183), .C(n1164), 
        .D(n1165), .Q(n1162) );
  XNR20 \i_iq_demod/filtre_Q/tot_adder/U45  ( .A(
        \i_iq_demod/filtre_Q/mult2 [5]), .B(\i_iq_demod/filtre_Q/mult1 [5]), 
        .Q(n1161) );
  OAI220 \i_iq_demod/filtre_Q/tot_adder/U44  ( .A(n233), .B(n188), .C(n1160), 
        .D(n1161), .Q(n1158) );
  XNR20 \i_iq_demod/filtre_Q/tot_adder/U40  ( .A(
        \i_iq_demod/filtre_Q/mult2 [7]), .B(\i_iq_demod/filtre_Q/mult1 [7]), 
        .Q(n1157) );
  OAI220 \i_iq_demod/filtre_Q/tot_adder/U39  ( .A(n232), .B(n187), .C(n1156), 
        .D(n1157), .Q(n1154) );
  XNR20 \i_iq_demod/filtre_Q/tot_adder/U35  ( .A(
        \i_iq_demod/filtre_Q/mult2 [9]), .B(\i_iq_demod/filtre_Q/mult1 [9]), 
        .Q(n1153) );
  OAI220 \i_iq_demod/filtre_Q/tot_adder/U34  ( .A(n1180), .B(n1181), .C(n1152), 
        .D(n1153), .Q(n1178) );
  XNR20 \i_iq_demod/filtre_Q/tot_adder/U29  ( .A(
        \i_iq_demod/filtre_Q/mult2 [11]), .B(\i_iq_demod/filtre_Q/mult1 [11]), 
        .Q(n1177) );
  XOR20 \i_iq_demod/filtre_Q/tot_adder/U28  ( .A(n1176), .B(n1177), .Q(
        \i_iq_demod/filtre_Q/tot [11]) );
  CLKIN0 \i_iq_demod/filtre_Q/tot_adder/U27  ( .A(
        \i_iq_demod/filtre_Q/mult2 [11]), .Q(n1174) );
  CLKIN0 \i_iq_demod/filtre_Q/tot_adder/U26  ( .A(
        \i_iq_demod/filtre_Q/mult1 [11]), .Q(n1175) );
  OAI220 \i_iq_demod/filtre_Q/tot_adder/U25  ( .A(n1174), .B(n1175), .C(n1176), 
        .D(n1177), .Q(n1171) );
  NOR20 \i_iq_demod/filtre_Q/tot_adder/U11  ( .A(n157), .B(n180), .Q(n1169) );
  XNR20 \i_iq_demod/filtre_Q/tot_adder/U10  ( .A(n1168), .B(n1169), .Q(
        \i_iq_demod/filtre_Q/tot [1]) );
  XOR20 \i_iq_demod/filtre_Q/tot_adder/U8  ( .A(n1164), .B(n1165), .Q(
        \i_iq_demod/filtre_Q/tot [3]) );
  XOR20 \i_iq_demod/filtre_Q/tot_adder/U6  ( .A(n1160), .B(n1161), .Q(
        \i_iq_demod/filtre_Q/tot [5]) );
  XOR20 \i_iq_demod/filtre_Q/tot_adder/U4  ( .A(n1156), .B(n1157), .Q(
        \i_iq_demod/filtre_Q/tot [7]) );
  XOR20 \i_iq_demod/filtre_Q/tot_adder/U2  ( .A(n1152), .B(n1153), .Q(
        \i_iq_demod/filtre_Q/tot [9]) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[12].adder/U39  ( .A(
        n1197), .B(\i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[12][0] ), .Q(\i_iq_demod/filtre_Q/mult2 [12]) );
  CLKIN0 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[12].adder/U37  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[12][0] ), .Q(n1149) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[12].adder/U36  ( .A(
        n1197), .B(n1149), .Q(n1151) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[11].adder/U39  ( .A(
        n1197), .B(\i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[11][0] ), .Q(\i_iq_demod/filtre_Q/mult2 [11]) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[11].adder/U38  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[11][1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[1] ), .Q(n1146) );
  CLKIN0 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[11].adder/U37  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[11][0] ), .Q(n1145) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[11].adder/U36  ( .A(
        n1197), .B(n1145), .Q(n1148) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[11].adder/U35  ( .A(
        n1146), .B(n1148), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[12][0] ) );
  NAND20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[11].adder/U34  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[11][1] ), .Q(n1147) );
  OAI310 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[11].adder/U33  ( .A(
        n1145), .B(n1146), .C(n1197), .D(n1147), .Q(n1143) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U39  ( .A(
        n1197), .B(\i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][0] ), .Q(\i_iq_demod/filtre_Q/mult2 [10]) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U38  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[1] ), .Q(n1140) );
  CLKIN0 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U37  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][0] ), .Q(n1139) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U36  ( .A(
        n1197), .B(n1139), .Q(n1142) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U35  ( .A(
        n1140), .B(n1142), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[11][0] ) );
  NAND20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U34  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][1] ), .Q(n1141) );
  OAI310 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U33  ( .A(
        n1139), .B(n1140), .C(n1197), .D(n1141), .Q(n1136) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U32  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[2] ), .Q(n1138) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U31  ( .A(
        n1136), .B(n1138), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[11][1] ) );
  CLKIN0 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U30  ( .A(
        n1138), .Q(n1137) );
  AOI220 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U29  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[2] ), .C(n1136), .D(
        n1137), .Q(n1134) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[10].adder/U28  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][3] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[3] ), .Q(n1135) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U39  ( .A(n1197), .B(\i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][0] ), .Q(
        \i_iq_demod/filtre_Q/mult2 [9]) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U38  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[1] ), .Q(n1131) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U36  ( .A(n1197), .B(n217), .Q(n1133) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U35  ( .A(n1131), .B(n1133), .Q(\i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][0] )
         );
  NAND20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U34  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][1] ), .Q(n1132)
         );
  OAI310 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U33  ( .A(n217), .B(n1131), .C(n1197), .D(n1132), .Q(n1128) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U32  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[2] ), .Q(n1130) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U31  ( .A(n1128), .B(n1130), .Q(\i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][1] )
         );
  CLKIN0 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U30  ( .A(
        n1130), .Q(n1129) );
  AOI220 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U29  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[2] ), .C(n1128), .D(
        n1129), .Q(n1126) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U28  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][3] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[3] ), .Q(n1127) );
  XOR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U27  ( .A(n1126), .B(n1127), .Q(\i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][2] )
         );
  OAI220 \i_iq_demod/filtre_Q/mult2_multiplier/genblk2[9].adder/U24  ( .A(n222), .B(n1195), .C(n1126), .D(n1127), .Q(n1125) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[8].adder/U39  ( .A(n1076), .B(\i_iq_demod/filtre_Q/mult2_multiplier/register[8][0] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [8]) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[8].adder/U36  ( .A(n1076), .B(n1121), .Q(n1124) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[8].adder/U35  ( .A(n1122), .B(n1124), .Q(\i_iq_demod/filtre_Q/mult2_multiplier/register[9][0] ) );
  NAND20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[8].adder/U34  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[8][1] ), .Q(n1123) );
  XOR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[8].adder/U27  ( .A(n1118), .B(n1746), .Q(\i_iq_demod/filtre_Q/mult2_multiplier/register[9][2] ) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[7].adder/U39  ( .A(n1076), .B(\i_iq_demod/filtre_Q/mult2_multiplier/register[7][0] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [7]) );
  CLKIN0 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[7].adder/U17  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[7][5] ), .Q(n1098) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[6].adder/U39  ( .A(n1076), .B(\i_iq_demod/filtre_Q/mult2_multiplier/register[6][0] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [6]) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[6].adder/U35  ( .A(n1094), .B(n1096), .Q(\i_iq_demod/filtre_Q/mult2_multiplier/register[7][0] ) );
  NAND20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[6].adder/U34  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[1] ), .B(n1779), .Q(
        n1095) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[5].adder/U39  ( .A(n1076), .B(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][0] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [5]) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[5].adder/U36  ( .A(n1076), .B(n1074), .Q(n1078) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[5].adder/U35  ( .A(n1075), .B(n1078), .Q(\i_iq_demod/filtre_Q/mult2_multiplier/register[6][0] ) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[4].adder/U39  ( .A(n1053), .B(\i_iq_demod/filtre_Q/mult2_multiplier/register[4][0] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [4]) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[3].adder/U39  ( .A(n1030), .B(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][0] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [3]) );
  CLKIN0 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[3].adder/U16  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[5] ), .Q(n1017) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[2].adder/U39  ( .A(n1008), .B(\i_iq_demod/filtre_Q/mult2_multiplier/register[2][0] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [2]) );
  CLKIN0 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[2].adder/U17  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][5] ), .Q(n993) );
  XNR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[1].adder/U39  ( .A(n1772), .B(\i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[1] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/S_pipe [1]) );
  NOR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[1].adder/U36  ( .A(n1772), .B(n981), .Q(n985) );
  CLKIN0 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[1].adder/U16  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[5] ), .Q(n970) );
  XOR20 \i_iq_demod/filtre_Q/mult2_multiplier/genblk1[1].adder/U10  ( .A(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[7] ), .Q(n966) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[12].adder/U39  ( .A(
        n1192), .B(\i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[12][0] ), .Q(\i_iq_demod/filtre_Q/mult1 [12]) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[12].adder/U37  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[12][0] ), .Q(n959)
         );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[12].adder/U36  ( .A(
        n1192), .B(n959), .Q(n961) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[11].adder/U39  ( .A(
        n1192), .B(\i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[11][0] ), .Q(\i_iq_demod/filtre_Q/mult1 [11]) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[11].adder/U37  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[11][0] ), .Q(n955)
         );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[11].adder/U36  ( .A(
        n1192), .B(n955), .Q(n958) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[11].adder/U35  ( .A(n956), .B(n958), .Q(\i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[12][0] ) );
  NAND20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[11].adder/U34  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[11][1] ), .Q(n957)
         );
  OAI310 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[11].adder/U33  ( .A(
        n955), .B(n956), .C(n1192), .D(n957), .Q(n953) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[10].adder/U39  ( .A(
        n1192), .B(\i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][0] ), .Q(\i_iq_demod/filtre_Q/mult1 [10]) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[10].adder/U37  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][0] ), .Q(n949)
         );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[10].adder/U36  ( .A(
        n1192), .B(n949), .Q(n952) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[10].adder/U35  ( .A(n950), .B(n952), .Q(\i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[11][0] ) );
  NAND20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[10].adder/U34  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][1] ), .Q(n951)
         );
  OAI310 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[10].adder/U33  ( .A(
        n949), .B(n950), .C(n1192), .D(n951), .Q(n946) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[10].adder/U32  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[2] ), .Q(n948) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[10].adder/U31  ( .A(n946), .B(n948), .Q(\i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[11][1] ) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[10].adder/U30  ( .A(
        n948), .Q(n947) );
  AOI220 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[10].adder/U29  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[2] ), .C(n946), .D(n947), .Q(n944) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[10].adder/U28  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][3] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[3] ), .Q(n945) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U39  ( .A(n1192), .B(\i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][0] ), .Q(
        \i_iq_demod/filtre_Q/mult1 [9]) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U38  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[1] ), .Q(n941) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U36  ( .A(n1192), .B(n216), .Q(n943) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U35  ( .A(n941), 
        .B(n943), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][0] ) );
  NAND20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U34  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][1] ), .Q(n942)
         );
  OAI310 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U33  ( .A(n216), .B(n941), .C(n1192), .D(n942), .Q(n938) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U32  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[2] ), .Q(n940) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U31  ( .A(n938), 
        .B(n940), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][1] ) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U30  ( .A(n940), .Q(n939) );
  AOI220 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U29  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[2] ), .C(n938), .D(n939), .Q(n936) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U28  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][3] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[3] ), .Q(n937) );
  XOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U27  ( .A(n936), 
        .B(n937), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][2] ) );
  OAI220 \i_iq_demod/filtre_Q/mult1_multiplier/genblk2[9].adder/U24  ( .A(n221), .B(n1189), .C(n936), .D(n937), .Q(n935) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[8].adder/U39  ( .A(n886), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/register[8][0] ), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [8]) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[8].adder/U36  ( .A(n886), 
        .B(n931), .Q(n934) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[8].adder/U35  ( .A(n932), 
        .B(n934), .Q(\i_iq_demod/filtre_Q/mult1_multiplier/register[9][0] ) );
  XOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[8].adder/U27  ( .A(n927), 
        .B(n928), .Q(\i_iq_demod/filtre_Q/mult1_multiplier/register[9][2] ) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[7].adder/U39  ( .A(n886), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/register[7][0] ), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [7]) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[7].adder/U36  ( .A(n886), 
        .B(n918), .Q(n921) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[7].adder/U35  ( .A(n919), 
        .B(n921), .Q(\i_iq_demod/filtre_Q/mult1_multiplier/register[8][0] ) );
  NAND20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[7].adder/U34  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[7][1] ), .Q(n920) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[6].adder/U39  ( .A(n886), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/register[6][0] ), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [6]) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[6].adder/U36  ( .A(n886), 
        .B(n903), .Q(n906) );
  NAND20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[6].adder/U34  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[6][1] ), .Q(n905) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[5].adder/U39  ( .A(n886), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/register[5][0] ), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [5]) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[5].adder/U36  ( .A(n886), 
        .B(n884), .Q(n888) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[5].adder/U16  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[5] ), .Q(n873) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[4].adder/U39  ( .A(n863), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][0] ), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [4]) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[4].adder/U16  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[5] ), .Q(n850) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[3].adder/U39  ( .A(n840), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/register[3][0] ), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [3]) );
  NOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[3].adder/U36  ( .A(n840), 
        .B(n838), .Q(n842) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[2].adder/U39  ( .A(n818), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][0] ), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [2]) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[2].adder/U26  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][3] ), .Q(n810) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[2].adder/U16  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[5] ), .Q(n805) );
  XNR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[1].adder/U39  ( .A(n1658), .B(\i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[1] ), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/S_pipe [1]) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[1].adder/U26  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[4] ), .Q(n786) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[1].adder/U25  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[3] ), .Q(n787) );
  CLKIN0 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[1].adder/U16  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[5] ), .Q(n781) );
  XOR20 \i_iq_demod/filtre_Q/mult1_multiplier/genblk1[1].adder/U10  ( .A(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[7] ), .Q(n777) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[12].adder/U39  ( .A(
        n1186), .B(\i_iq_demod/filtre_I/mult2_multiplier/register_pipe[12][0] ), .Q(\i_iq_demod/filtre_I/mult2 [12]) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[12].adder/U37  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[12][0] ), .Q(n770)
         );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[12].adder/U36  ( .A(
        n1186), .B(n770), .Q(n772) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[11].adder/U39  ( .A(
        n1186), .B(\i_iq_demod/filtre_I/mult2_multiplier/register_pipe[11][0] ), .Q(\i_iq_demod/filtre_I/mult2 [11]) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[11].adder/U38  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[11][1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[1] ), .Q(n767) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[11].adder/U37  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[11][0] ), .Q(n766)
         );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[11].adder/U36  ( .A(
        n1186), .B(n766), .Q(n769) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[11].adder/U35  ( .A(n767), .B(n769), .Q(\i_iq_demod/filtre_I/mult2_multiplier/register_pipe[12][0] ) );
  NAND20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[11].adder/U34  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[11][1] ), .Q(n768)
         );
  OAI310 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[11].adder/U33  ( .A(
        n766), .B(n767), .C(n1186), .D(n768), .Q(n764) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U39  ( .A(
        n1186), .B(\i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][0] ), .Q(\i_iq_demod/filtre_I/mult2 [10]) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U38  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[1] ), .Q(n761) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U37  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][0] ), .Q(n760)
         );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U36  ( .A(
        n1186), .B(n760), .Q(n763) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U35  ( .A(n761), .B(n763), .Q(\i_iq_demod/filtre_I/mult2_multiplier/register_pipe[11][0] ) );
  NAND20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U34  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][1] ), .Q(n762)
         );
  OAI310 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U33  ( .A(
        n760), .B(n761), .C(n1186), .D(n762), .Q(n757) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U32  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[2] ), .Q(n759) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U31  ( .A(n757), .B(n759), .Q(\i_iq_demod/filtre_I/mult2_multiplier/register_pipe[11][1] ) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U30  ( .A(
        n759), .Q(n758) );
  AOI220 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U29  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[2] ), .C(n757), .D(n758), .Q(n755) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[10].adder/U28  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][3] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[3] ), .Q(n756) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U39  ( .A(n1186), .B(\i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][0] ), .Q(
        \i_iq_demod/filtre_I/mult2 [9]) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U38  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[1] ), .Q(n752) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U36  ( .A(n1186), .B(n215), .Q(n754) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U35  ( .A(n752), 
        .B(n754), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][0] ) );
  NAND20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U34  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][1] ), .Q(n753)
         );
  OAI310 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U33  ( .A(n215), .B(n752), .C(n1186), .D(n753), .Q(n749) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U32  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[2] ), .Q(n751) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U31  ( .A(n749), 
        .B(n751), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][1] ) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U30  ( .A(n751), .Q(n750) );
  AOI220 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U29  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[2] ), .C(n749), .D(n750), .Q(n747) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U28  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][3] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[3] ), .Q(n748) );
  XOR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U27  ( .A(n747), 
        .B(n748), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][2] ) );
  OAI220 \i_iq_demod/filtre_I/mult2_multiplier/genblk2[9].adder/U24  ( .A(n220), .B(n1184), .C(n747), .D(n748), .Q(n746) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[8].adder/U39  ( .A(n697), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/register[8][0] ), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [8]) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[8].adder/U35  ( .A(n743), 
        .B(n745), .Q(\i_iq_demod/filtre_I/mult2_multiplier/register[9][0] ) );
  XOR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[8].adder/U27  ( .A(n1631), .B(n1623), .Q(\i_iq_demod/filtre_I/mult2_multiplier/register[9][2] ) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[7].adder/U39  ( .A(n697), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/register[7][0] ), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [7]) );
  NOR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[7].adder/U36  ( .A(n697), 
        .B(n729), .Q(n732) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[7].adder/U35  ( .A(n730), 
        .B(n732), .Q(\i_iq_demod/filtre_I/mult2_multiplier/register[8][0] ) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[7].adder/U17  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register[7][5] ), .Q(n719) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[6].adder/U39  ( .A(n697), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/register[6][0] ), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [6]) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[5].adder/U39  ( .A(n697), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/register[5][0] ), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [5]) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[5].adder/U35  ( .A(n696), 
        .B(n699), .Q(\i_iq_demod/filtre_I/mult2_multiplier/register[6][0] ) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[4].adder/U39  ( .A(n674), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/register[4][0] ), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [4]) );
  NAND20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[4].adder/U34  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][1] ), .Q(n675) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[3].adder/U35  ( .A(n650), 
        .B(n653), .Q(\i_iq_demod/filtre_I/mult2_multiplier/register[4][0] ) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[2].adder/U39  ( .A(n629), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/register[2][0] ), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [2]) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[2].adder/U26  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][3] ), .Q(n621) );
  XNR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[1].adder/U39  ( .A(n1715), .B(\i_iq_demod/filtre_I/mult2_multiplier/_0_net_[1] ), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/S_pipe [1]) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[1].adder/U26  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[4] ), .Q(n596) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[1].adder/U25  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[3] ), .Q(n597) );
  CLKIN0 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[1].adder/U16  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[5] ), .Q(n591) );
  XOR20 \i_iq_demod/filtre_I/mult2_multiplier/genblk1[1].adder/U10  ( .A(
        \i_iq_demod/filtre_I/mult2_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[7] ), .Q(n587) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[12].adder/U39  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/n21 ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[12][0] ), .Q(
        \i_iq_demod/filtre_I/mult1 [12]) );
  CLKIN0 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[12].adder/U37  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[12][0] ), .Q(n580)
         );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[12].adder/U36  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/n21 ), .B(n580), .Q(n582) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[11].adder/U39  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/n21 ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[11][0] ), .Q(
        \i_iq_demod/filtre_I/mult1 [11]) );
  CLKIN0 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[11].adder/U37  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[11][0] ), .Q(n576)
         );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[11].adder/U36  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/n21 ), .B(n576), .Q(n579) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[11].adder/U35  ( .A(n577), .B(n579), .Q(\i_iq_demod/filtre_I/mult1_multiplier/register_pipe[12][0] ) );
  NAND20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[11].adder/U34  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[11][1] ), .Q(n578)
         );
  OAI310 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[11].adder/U33  ( .A(
        n576), .B(n577), .C(\i_iq_demod/filtre_I/mult1_multiplier/n21 ), .D(
        n578), .Q(n574) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[10].adder/U39  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/n21 ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][0] ), .Q(
        \i_iq_demod/filtre_I/mult1 [10]) );
  CLKIN0 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[10].adder/U37  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][0] ), .Q(n570)
         );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[10].adder/U36  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/n21 ), .B(n570), .Q(n573) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[10].adder/U35  ( .A(n571), .B(n573), .Q(\i_iq_demod/filtre_I/mult1_multiplier/register_pipe[11][0] ) );
  NAND20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[10].adder/U34  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][1] ), .Q(n572)
         );
  OAI310 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[10].adder/U33  ( .A(
        n570), .B(n571), .C(\i_iq_demod/filtre_I/mult1_multiplier/n21 ), .D(
        n572), .Q(n567) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[10].adder/U32  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[2] ), .Q(n569) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[10].adder/U31  ( .A(n567), .B(n569), .Q(\i_iq_demod/filtre_I/mult1_multiplier/register_pipe[11][1] ) );
  CLKIN0 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[10].adder/U30  ( .A(
        n569), .Q(n568) );
  AOI220 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[10].adder/U29  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[2] ), .C(n567), .D(n568), .Q(n565) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[10].adder/U28  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][3] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[3] ), .Q(n566) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U39  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/n21 ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][0] ), .Q(
        \i_iq_demod/filtre_I/mult1 [9]) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U38  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[1] ), .Q(n562) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U36  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/n21 ), .B(n214), .Q(n564) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U35  ( .A(n562), 
        .B(n564), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][0] ) );
  NAND20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U34  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][1] ), .Q(n563)
         );
  OAI310 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U33  ( .A(n214), .B(n562), .C(\i_iq_demod/filtre_I/mult1_multiplier/n21 ), .D(n563), .Q(n559)
         );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U32  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[2] ), .Q(n561) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U31  ( .A(n559), 
        .B(n561), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][1] ) );
  CLKIN0 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U30  ( .A(n561), .Q(n560) );
  AOI220 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U29  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[2] ), .C(n559), .D(n560), .Q(n557) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U28  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][3] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[3] ), .Q(n558) );
  XOR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U27  ( .A(n557), 
        .B(n558), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][2] ) );
  OAI220 \i_iq_demod/filtre_I/mult1_multiplier/genblk2[9].adder/U24  ( .A(n219), .B(\i_iq_demod/filtre_I/mult1_multiplier/n18 ), .C(n557), .D(n558), .Q(n556)
         );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[8].adder/U39  ( .A(n507), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/register[8][0] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [8]) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[8].adder/U36  ( .A(n507), 
        .B(n552), .Q(n555) );
  NAND20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[8].adder/U34  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[1] ), .B(n1717), .Q(
        n554) );
  XOR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[8].adder/U27  ( .A(n1723), .B(n549), .Q(\i_iq_demod/filtre_I/mult1_multiplier/register[9][2] ) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[7].adder/U39  ( .A(n507), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/register[7][0] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [7]) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[7].adder/U36  ( .A(n507), 
        .B(n539), .Q(n542) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[7].adder/U35  ( .A(n540), 
        .B(n542), .Q(\i_iq_demod/filtre_I/mult1_multiplier/register[8][0] ) );
  NAND20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[7].adder/U34  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[7][1] ), .Q(n541) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[6].adder/U39  ( .A(n507), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/register[6][0] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [6]) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[6].adder/U35  ( .A(n525), 
        .B(n527), .Q(\i_iq_demod/filtre_I/mult1_multiplier/register[7][0] ) );
  NAND20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[6].adder/U34  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[6][1] ), .Q(n526) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[5].adder/U39  ( .A(n507), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/register[5][0] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [5]) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[5].adder/U36  ( .A(n507), 
        .B(n505), .Q(n509) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[4].adder/U39  ( .A(n484), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/register[4][0] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [4]) );
  CLKIN0 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[4].adder/U16  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[5] ), .Q(n471) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[3].adder/U39  ( .A(n461), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/register[3][0] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [3]) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[3].adder/U35  ( .A(n460), 
        .B(n463), .Q(\i_iq_demod/filtre_I/mult1_multiplier/register[4][0] ) );
  NAND20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[3].adder/U34  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][1] ), .Q(n462) );
  CLKIN0 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[3].adder/U17  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][5] ), .Q(n447) );
  CLKIN0 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[3].adder/U16  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[5] ), .Q(n448) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[1].adder/U39  ( .A(n415), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/_0_net_[1] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [1]) );
  CLKIN0 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[1].adder/U16  ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[5] ), .Q(n402) );
  ADD22 \i_cdr/i_cdr/add_119/U1_1_1  ( .A(\i_cdr/i_cdr/count [1]), .B(
        \i_cdr/i_cdr/count [0]), .CO(\i_cdr/i_cdr/add_119/carry [2]), .S(
        \i_cdr/i_cdr/N149 ) );
  ADD22 \i_cdr/i_cdr/add_119/U1_1_2  ( .A(\i_cdr/i_cdr/count [2]), .B(
        \i_cdr/i_cdr/add_119/carry [2]), .CO(\i_cdr/i_cdr/add_119/carry [3]), 
        .S(\i_cdr/i_cdr/N150 ) );
  ADD22 \i_cdr/i_cdr/add_119/U1_1_3  ( .A(\i_cdr/i_cdr/count [3]), .B(
        \i_cdr/i_cdr/add_119/carry [3]), .CO(\i_cdr/i_cdr/add_119/carry [4]), 
        .S(\i_cdr/i_cdr/N151 ) );
  ADD32 \i_cordic/S1/sub_50/U2_2  ( .A(\i_cordic/cor_x_s0[1][2] ), .B(
        \i_cordic/S1/sub_50/B_not [2]), .CI(\i_cordic/S1/sub_50/carry [2]), 
        .CO(\i_cordic/S1/sub_50/carry [3]), .S(\i_cordic/S1/N11 ) );
  ADD32 \i_cordic/S1/sub_50/U2_3  ( .A(\i_cordic/cor_x_s0[1][3] ), .B(
        \i_cordic/S1/sub_50/B_not [3]), .CI(\i_cordic/S1/sub_50/carry [3]), 
        .CO(\i_cordic/S1/sub_50/carry [4]), .S(\i_cordic/S1/N12 ) );
  ADD32 \i_cordic/S1/sub_50/U2_4  ( .A(\i_cordic/cor_x_s0[1][4] ), .B(
        \i_cordic/S1/sub_50/B_not [5]), .CI(\i_cordic/S1/sub_50/carry [4]), 
        .CO(\i_cordic/S1/sub_50/carry [5]), .S(\i_cordic/S1/N13 ) );
  ADD32 \i_cordic/S1/sub_53/U2_1  ( .A(\i_cordic/cor_y_s0[1][1] ), .B(
        \i_cordic/S1/sub_53/B_not [1]), .CI(\i_cordic/S1/sub_53/carry [1]), 
        .CO(\i_cordic/S1/sub_53/carry [2]), .S(\i_cordic/S1/N16 ) );
  ADD32 \i_cordic/S1/sub_53/U2_2  ( .A(\i_cordic/cor_y_s0[1][2] ), .B(
        \i_cordic/S1/sub_53/B_not [2]), .CI(\i_cordic/S1/sub_53/carry [2]), 
        .CO(\i_cordic/S1/sub_53/carry [3]), .S(\i_cordic/S1/N17 ) );
  ADD32 \i_cordic/S1/sub_53/U2_3  ( .A(\i_cordic/cor_y_s0[1][3] ), .B(
        \i_cordic/S1/sub_53/B_not [3]), .CI(\i_cordic/S1/sub_53/carry [3]), 
        .CO(\i_cordic/S1/sub_53/carry [4]), .S(\i_cordic/S1/N18 ) );
  ADD32 \i_cordic/S1/sub_53/U2_4  ( .A(\i_cordic/cor_y_s0[1][4] ), .B(
        \i_cordic/S1/sub_53/B_not [5]), .CI(\i_cordic/S1/sub_53/carry [4]), 
        .CO(\i_cordic/S1/sub_53/carry [5]), .S(\i_cordic/S1/N19 ) );
  ADD32 \i_cordic/S0/r64/U1_1  ( .A(\i_cordic/cor_x_s0[0][1] ), .B(
        \i_cordic/cor_y_s0[0][1] ), .CI(\i_cordic/S0/r64/carry [1]), .CO(
        \i_cordic/S0/r64/carry [2]), .S(\i_cordic/S0/N4 ) );
  ADD32 \i_cordic/S0/r64/U1_2  ( .A(\i_cordic/cor_x_s0[0][2] ), .B(
        \i_cordic/cor_y_s0[0][2] ), .CI(\i_cordic/S0/r64/carry [2]), .CO(
        \i_cordic/S0/r64/carry [3]), .S(\i_cordic/S0/N5 ) );
  ADD32 \i_cordic/S0/r64/U1_3  ( .A(\i_cordic/cor_x_s0[0][3] ), .B(
        \i_cordic/cor_y_s0[0][3] ), .CI(\i_cordic/S0/r64/carry [3]), .CO(
        \i_cordic/S0/r64/carry [4]), .S(\i_cordic/S0/N6 ) );
  ADD32 \i_cordic/S0/r64/U1_4  ( .A(n275), .B(\i_cordic/cor_y_s0[0][4] ), .CI(
        \i_cordic/S0/r64/carry [4]), .CO(\i_cordic/S0/r64/carry [5]), .S(
        \i_cordic/S0/N7 ) );
  ADD32 \i_cordic/S0/sub_50/U2_1  ( .A(\i_cordic/cor_x_s0[0][1] ), .B(
        \i_cordic/S0/sub_50/B_not [1]), .CI(\i_cordic/S0/sub_50/carry [1]), 
        .CO(\i_cordic/S0/sub_50/carry [2]), .S(\i_cordic/S0/N10 ) );
  ADD32 \i_cordic/S0/sub_50/U2_2  ( .A(\i_cordic/cor_x_s0[0][2] ), .B(
        \i_cordic/S0/sub_50/B_not [2]), .CI(\i_cordic/S0/sub_50/carry [2]), 
        .CO(\i_cordic/S0/sub_50/carry [3]), .S(\i_cordic/S0/N11 ) );
  ADD32 \i_cordic/S0/sub_50/U2_3  ( .A(\i_cordic/cor_x_s0[0][3] ), .B(
        \i_cordic/S0/sub_50/B_not [3]), .CI(\i_cordic/S0/sub_50/carry [3]), 
        .CO(\i_cordic/S0/sub_50/carry [4]), .S(\i_cordic/S0/N12 ) );
  ADD32 \i_cordic/S0/sub_50/U2_4  ( .A(n275), .B(\i_cordic/S0/sub_50/B_not [4]), .CI(\i_cordic/S0/sub_50/carry [4]), .CO(\i_cordic/S0/sub_50/carry [5]), .S(
        \i_cordic/S0/N13 ) );
  ADD32 \i_cordic/S0/sub_53/U2_1  ( .A(\i_cordic/cor_y_s0[0][1] ), .B(
        \i_cordic/n21 ), .CI(\i_cordic/S0/sub_53/carry [1]), .CO(
        \i_cordic/S0/sub_53/carry [2]), .S(\i_cordic/S0/N16 ) );
  ADD32 \i_cordic/S0/sub_53/U2_2  ( .A(\i_cordic/cor_y_s0[0][2] ), .B(
        \i_cordic/n20 ), .CI(\i_cordic/S0/sub_53/carry [2]), .CO(
        \i_cordic/S0/sub_53/carry [3]), .S(\i_cordic/S0/N17 ) );
  ADD32 \i_cordic/S0/sub_53/U2_3  ( .A(\i_cordic/cor_y_s0[0][3] ), .B(
        \i_cordic/n19 ), .CI(\i_cordic/S0/sub_53/carry [3]), .CO(
        \i_cordic/S0/sub_53/carry [4]), .S(\i_cordic/S0/N18 ) );
  ADD32 \i_cordic/S0/sub_53/U2_4  ( .A(\i_cordic/cor_y_s0[0][4] ), .B(n89), 
        .CI(\i_cordic/S0/sub_53/carry [4]), .CO(\i_cordic/S0/sub_53/carry [5]), 
        .S(\i_cordic/S0/N19 ) );
  ADD32 \i_iq_demod/demod/dp_cluster_0/sub_88/U2_1  ( .A(
        \i_iq_demod/demod/QC [1]), .B(
        \i_iq_demod/demod/dp_cluster_0/sub_88/B_not [1]), .CI(
        \i_iq_demod/demod/dp_cluster_0/sub_88/carry [1]), .CO(
        \i_iq_demod/demod/dp_cluster_0/sub_88/carry [2]), .S(
        \i_iq_demod/demod/dp_cluster_0/N90 ) );
  ADD32 \i_iq_demod/demod/dp_cluster_0/sub_88/U2_2  ( .A(
        \i_iq_demod/demod/QC [2]), .B(
        \i_iq_demod/demod/dp_cluster_0/sub_88/B_not [2]), .CI(
        \i_iq_demod/demod/dp_cluster_0/sub_88/carry [2]), .CO(
        \i_iq_demod/demod/dp_cluster_0/sub_88/carry [3]), .S(
        \i_iq_demod/demod/dp_cluster_0/N91 ) );
  ADD32 \i_iq_demod/demod/dp_cluster_0/sub_88/U2_3  ( .A(
        \i_iq_demod/demod/QC [3]), .B(
        \i_iq_demod/demod/dp_cluster_0/sub_88/B_not [3]), .CI(
        \i_iq_demod/demod/dp_cluster_0/sub_88/carry [3]), .CO(
        \i_iq_demod/demod/dp_cluster_0/sub_88/carry [4]), .S(
        \i_iq_demod/demod/dp_cluster_0/N92 ) );
  ADD32 \i_iq_demod/demod/dp_cluster_0/sub_88/U2_4  ( .A(
        \i_iq_demod/demod/QC [4]), .B(
        \i_iq_demod/demod/dp_cluster_0/sub_88/B_not [4]), .CI(
        \i_iq_demod/demod/dp_cluster_0/sub_88/carry [4]), .S(
        \i_iq_demod/demod/dp_cluster_0/N93 ) );
  ADD32 \i_iq_demod/demod/dp_cluster_1/add_87/U1_1  ( .A(
        \i_iq_demod/demod/IC [1]), .B(\i_iq_demod/demod/QS [1]), .CI(
        \i_iq_demod/demod/dp_cluster_1/add_87/carry [1]), .CO(
        \i_iq_demod/demod/dp_cluster_1/add_87/carry [2]), .S(
        \i_iq_demod/demod/dp_cluster_1/N85 ) );
  ADD32 \i_iq_demod/demod/dp_cluster_1/add_87/U1_2  ( .A(
        \i_iq_demod/demod/IC [2]), .B(\i_iq_demod/demod/QS [2]), .CI(
        \i_iq_demod/demod/dp_cluster_1/add_87/carry [2]), .CO(
        \i_iq_demod/demod/dp_cluster_1/add_87/carry [3]), .S(
        \i_iq_demod/demod/dp_cluster_1/N86 ) );
  ADD32 \i_iq_demod/demod/dp_cluster_1/add_87/U1_3  ( .A(
        \i_iq_demod/demod/IC [3]), .B(\i_iq_demod/demod/QS [3]), .CI(
        \i_iq_demod/demod/dp_cluster_1/add_87/carry [3]), .CO(
        \i_iq_demod/demod/dp_cluster_1/add_87/carry [4]), .S(
        \i_iq_demod/demod/dp_cluster_1/N87 ) );
  ADD32 \i_iq_demod/demod/dp_cluster_1/add_87/U1_4  ( .A(
        \i_iq_demod/demod/IC [4]), .B(\i_iq_demod/demod/QS [4]), .CI(
        \i_iq_demod/demod/dp_cluster_1/add_87/carry [4]), .S(
        \i_iq_demod/demod/dp_cluster_1/N88 ) );
  ADD22 \i_fifo_rx/add_90/U1_1_1  ( .A(\i_fifo_rx/i [1]), .B(\i_fifo_rx/i [0]), 
        .CO(\i_fifo_rx/add_90/carry [2]), .S(\i_fifo_rx/N54 ) );
  ADD22 \i_fifo_rx/add_90/U1_1_2  ( .A(\i_fifo_rx/i [2]), .B(
        \i_fifo_rx/add_90/carry [2]), .CO(\i_fifo_rx/add_90/carry [3]), .S(
        \i_fifo_rx/N55 ) );
  ADD22 \i_fifo_rx/add_90/U1_1_3  ( .A(\i_fifo_rx/i [3]), .B(
        \i_fifo_rx/add_90/carry [3]), .CO(\i_fifo_rx/add_90/carry [4]), .S(
        \i_fifo_rx/N56 ) );
  ADD22 \i_fifo_rx/add_90/U1_1_4  ( .A(\i_fifo_rx/i [4]), .B(
        \i_fifo_rx/add_90/carry [4]), .CO(\i_fifo_rx/add_90/carry [5]), .S(
        \i_fifo_rx/N57 ) );
  ADD22 \i_fifo_rx/add_90/U1_1_5  ( .A(\i_fifo_rx/i [5]), .B(
        \i_fifo_rx/add_90/carry [5]), .CO(\i_fifo_rx/add_90/carry [6]), .S(
        \i_fifo_rx/N58 ) );
  ADD22 \i_fifo_rx/add_90/U1_1_6  ( .A(\i_fifo_rx/i [6]), .B(
        \i_fifo_rx/add_90/carry [6]), .CO(\i_fifo_rx/add_90/carry [7]), .S(
        \i_fifo_rx/N59 ) );
  ADD22 \i_fifo_rx/add_106/U1_1_1  ( .A(n305), .B(n302), .CO(
        \i_fifo_rx/add_106/carry [2]), .S(\i_fifo_rx/N81 ) );
  ADD22 \i_fifo_rx/add_106/U1_1_3  ( .A(n274), .B(\i_fifo_rx/add_106/carry [3]), .CO(\i_fifo_rx/add_106/carry [4]), .S(\i_fifo_rx/N83 ) );
  ADD22 \i_fifo_rx/add_106/U1_1_4  ( .A(\i_fifo_rx/N37 ), .B(
        \i_fifo_rx/add_106/carry [4]), .CO(\i_fifo_rx/add_106/carry [5]), .S(
        \i_fifo_rx/N84 ) );
  ADD22 \i_fifo_rx/add_106/U1_1_5  ( .A(\i_fifo_rx/N38 ), .B(
        \i_fifo_rx/add_106/carry [5]), .CO(\i_fifo_rx/add_106/carry [6]), .S(
        \i_fifo_rx/N85 ) );
  ADD22 \i_fifo_rx/add_139/U1_1_1  ( .A(n311), .B(\i_fifo_rx/N39 ), .CO(
        \i_fifo_rx/add_139/carry [2]), .S(\i_fifo_rx/N689 ) );
  ADD22 \i_fifo_rx/add_139/U1_1_2  ( .A(\i_fifo_rx/N41 ), .B(
        \i_fifo_rx/add_139/carry [2]), .CO(\i_fifo_rx/add_139/carry [3]), .S(
        \i_fifo_rx/N690 ) );
  ADD22 \i_fifo_rx/add_139/U1_1_5  ( .A(\i_fifo_rx/N44 ), .B(
        \i_fifo_rx/add_139/carry [5]), .CO(\i_fifo_rx/add_139/carry [6]), .S(
        \i_fifo_rx/N693 ) );
  ADD22 \i_fifo_tx/r80/U1_1_1  ( .A(\i_fifo_tx/counter_clock [1]), .B(
        \i_fifo_tx/counter_clock [0]), .CO(\i_fifo_tx/r80/carry [2]), .S(
        \i_fifo_tx/N149 ) );
  ADD22 \i_fifo_tx/r80/U1_1_2  ( .A(\i_fifo_tx/counter_clock [2]), .B(
        \i_fifo_tx/r80/carry [2]), .CO(\i_fifo_tx/r80/carry [3]), .S(
        \i_fifo_tx/N150 ) );
  ADD22 \i_fifo_tx/r80/U1_1_3  ( .A(\i_fifo_tx/counter_clock [3]), .B(
        \i_fifo_tx/r80/carry [3]), .CO(\i_fifo_tx/r80/carry [4]), .S(
        \i_fifo_tx/N151 ) );
  ADD22 \i_fifo_tx/add_100/U1_1_1  ( .A(n318), .B(n317), .CO(
        \i_fifo_tx/add_100/carry [2]), .S(\i_fifo_tx/N129 ) );
  ADD22 \i_fifo_tx/add_100/U1_1_3  ( .A(n273), .B(\i_fifo_tx/add_100/carry [3]), .CO(\i_fifo_tx/add_100/carry [4]), .S(\i_fifo_tx/N131 ) );
  ADD22 \i_fifo_tx/add_100/U1_1_4  ( .A(\i_fifo_tx/N28 ), .B(
        \i_fifo_tx/add_100/carry [4]), .CO(\i_fifo_tx/add_100/carry [5]), .S(
        \i_fifo_tx/N132 ) );
  ADD22 \i_fifo_tx/add_100/U1_1_5  ( .A(\i_fifo_tx/N29 ), .B(
        \i_fifo_tx/add_100/carry [5]), .CO(\i_fifo_tx/add_100/carry [6]), .S(
        \i_fifo_tx/N133 ) );
  ADD22 \i_fifo_tx/add_180/U1_1_1  ( .A(n328), .B(\i_fifo_tx/N30 ), .CO(
        \i_fifo_tx/add_180/carry [2]), .S(\i_fifo_tx/N156 ) );
  ADD22 \i_fifo_tx/add_180/U1_1_4  ( .A(\i_fifo_tx/N34 ), .B(
        \i_fifo_tx/add_180/carry [4]), .CO(\i_fifo_tx/add_180/carry [5]), .S(
        \i_fifo_tx/N159 ) );
  ADD22 \i_fifo_tx/add_180/U1_1_5  ( .A(\i_fifo_tx/N35 ), .B(
        \i_fifo_tx/add_180/carry [5]), .CO(\i_fifo_tx/add_180/carry [6]), .S(
        \i_fifo_tx/N160 ) );
  DFEC1 \i_fifo_tx/wr_ptr_reg[6]  ( .D(\i_fifo_tx/N134 ), .E(\i_fifo_tx/n152 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/wr_ptr[6] ), .QN(
        \i_fifo_tx/n183 ) );
  DFEC1 \i_fifo_tx/rd_ptr_reg[6]  ( .D(\i_fifo_tx/N161 ), .E(\i_fifo_tx/n187 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/rd_ptr[6] ), .QN(
        \i_fifo_tx/n188 ) );
  DFEC1 \i_fifo_rx/mem_reg[0][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n168 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[0][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[1][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n166 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[1][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[2][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n164 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[2][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[3][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n162 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[3][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[4][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n160 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[4][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[5][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n158 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[5][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[6][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n156 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[6][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[7][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n150 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[7][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[8][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n148 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[8][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[9][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n146 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[9][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[10][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n144 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[10][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[11][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n142 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[11][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[12][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n140 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[12][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[13][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n138 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[13][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[14][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n136 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[14][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[15][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n133 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[15][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[16][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n131 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[16][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[17][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n129 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[17][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[18][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n127 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[18][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[19][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n125 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[19][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[20][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n123 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[20][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[21][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n121 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[21][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[22][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n119 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[22][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[23][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n116 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[23][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[25][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n112 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[25][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[26][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n110 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[26][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[27][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n108 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[27][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[28][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n106 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[28][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[29][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n104 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[29][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[30][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n102 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[30][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[31][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n99 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[31][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[32][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n97 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[32][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[33][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n95 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[33][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[34][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n93 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[34][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[35][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[35][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[36][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n89 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[36][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[37][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n87 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[37][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[38][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n85 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[38][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[39][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n82 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[39][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[40][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n80 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[40][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[41][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n78 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[41][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[42][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n76 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[42][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[43][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[43][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[44][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[44][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[45][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[45][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[46][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[46][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[47][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[47][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[48][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[48][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[49][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[49][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[50][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[50][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[51][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[51][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[52][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[52][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[53][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[53][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[54][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[54][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[55][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[55][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[56][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[56][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[57][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[57][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[58][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[58][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[59][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[59][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[60][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[60][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[61][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[61][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[62][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[62][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[63][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[63][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[24][0]  ( .D(\i_fifo_rx/n3 ), .E(\i_fifo_rx/n114 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[24][0] ) );
  DFEC1 \i_fifo_rx/mem_reg[0][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n168 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[0][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[1][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n166 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[1][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[2][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n164 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[2][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[3][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n162 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[3][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[4][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n160 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[4][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[5][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n158 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[5][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[6][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n156 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[6][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[7][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n150 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[7][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[8][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n148 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[8][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[9][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n146 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[9][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[10][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n144 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[10][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[11][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n142 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[11][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[12][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n140 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[12][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[13][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n138 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[13][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[14][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n136 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[14][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[15][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n133 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[15][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[16][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n131 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[16][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[17][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n129 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[17][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[18][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n127 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[18][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[19][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n125 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[19][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[20][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n123 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[20][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[21][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n121 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[21][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[22][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n119 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[22][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[23][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n116 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[23][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[25][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n112 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[25][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[26][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n110 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[26][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[27][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n108 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[27][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[28][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n106 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[28][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[29][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n104 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[29][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[30][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n102 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[30][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[31][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n99 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[31][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[32][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n97 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[32][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[33][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n95 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[33][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[34][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n93 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[34][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[35][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[35][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[36][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n89 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[36][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[37][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n87 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[37][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[38][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n85 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[38][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[39][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n82 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[39][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[40][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n80 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[40][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[41][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n78 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[41][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[42][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n76 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[42][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[43][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[43][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[44][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[44][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[45][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[45][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[46][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[46][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[47][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[47][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[48][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[48][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[49][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[49][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[50][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[50][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[51][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[51][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[52][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[52][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[53][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[53][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[54][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[54][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[55][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[55][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[56][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[56][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[57][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[57][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[58][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[58][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[59][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[59][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[60][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[60][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[61][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[61][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[62][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[62][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[63][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[63][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[24][1]  ( .D(\i_fifo_rx/n4 ), .E(\i_fifo_rx/n114 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[24][1] ) );
  DFEC1 \i_fifo_rx/mem_reg[0][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n168 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[0][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[1][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n166 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[1][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[2][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n164 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[2][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[3][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n162 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[3][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[4][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n160 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[4][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[5][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n158 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[5][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[6][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n156 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[6][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[7][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n150 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[7][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[8][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n148 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[8][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[9][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n146 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[9][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[10][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n144 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[10][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[11][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n142 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[11][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[12][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n140 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[12][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[13][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n138 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[13][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[14][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n136 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[14][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[15][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n133 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[15][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[16][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n131 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[16][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[17][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n129 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[17][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[18][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n127 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[18][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[19][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n125 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[19][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[20][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n123 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[20][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[21][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n121 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[21][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[22][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n119 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[22][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[23][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n116 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[23][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[25][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n112 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[25][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[26][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n110 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[26][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[27][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n108 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[27][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[28][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n106 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[28][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[29][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n104 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[29][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[30][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n102 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[30][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[31][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n99 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[31][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[32][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n97 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[32][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[33][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n95 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[33][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[34][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n93 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[34][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[35][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[35][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[36][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n89 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[36][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[37][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n87 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[37][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[38][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n85 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[38][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[39][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n82 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[39][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[40][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n80 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[40][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[41][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n78 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[41][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[42][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n76 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[42][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[43][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[43][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[44][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[44][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[45][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[45][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[46][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[46][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[47][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[47][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[48][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[48][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[49][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[49][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[50][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[50][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[51][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[51][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[52][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[52][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[53][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[53][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[54][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[54][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[55][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[55][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[56][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[56][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[57][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[57][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[58][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[58][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[59][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[59][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[60][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[60][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[61][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[61][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[62][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[62][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[63][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[63][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[24][2]  ( .D(\i_fifo_rx/n5 ), .E(\i_fifo_rx/n114 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[24][2] ) );
  DFEC1 \i_fifo_rx/mem_reg[0][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n168 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[0][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[1][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n166 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[1][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[2][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n164 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[2][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[3][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n162 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[3][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[4][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n160 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[4][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[5][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n158 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[5][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[6][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n156 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[6][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[7][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n150 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[7][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[8][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n148 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[8][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[9][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n146 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[9][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[10][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n144 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[10][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[11][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n142 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[11][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[12][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n140 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[12][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[13][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n138 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[13][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[14][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n136 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[14][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[15][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n133 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[15][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[16][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n131 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[16][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[17][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n129 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[17][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[18][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n127 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[18][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[19][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n125 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[19][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[20][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n123 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[20][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[21][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n121 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[21][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[22][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n119 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[22][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[23][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n116 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[23][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[25][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n112 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[25][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[26][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n110 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[26][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[27][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n108 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[27][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[28][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n106 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[28][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[29][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n104 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[29][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[30][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n102 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[30][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[31][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n99 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[31][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[32][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n97 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[32][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[33][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n95 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[33][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[34][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n93 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[34][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[35][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[35][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[36][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n89 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[36][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[37][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n87 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[37][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[38][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n85 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[38][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[39][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n82 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[39][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[40][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n80 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[40][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[41][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n78 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[41][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[42][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n76 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[42][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[43][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[43][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[44][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[44][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[45][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[45][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[46][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[46][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[47][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[47][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[48][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[48][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[49][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[49][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[50][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[50][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[51][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[51][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[52][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[52][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[53][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[53][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[54][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[54][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[55][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[55][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[56][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[56][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[57][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[57][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[58][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[58][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[59][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[59][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[60][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[60][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[61][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[61][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[62][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[62][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[63][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[63][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[24][3]  ( .D(\i_fifo_rx/n6 ), .E(\i_fifo_rx/n114 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[24][3] ) );
  DFEC1 \i_fifo_rx/mem_reg[0][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n168 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[0][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[1][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n166 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[1][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[2][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n164 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[2][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[3][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n162 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[3][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[4][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n160 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[4][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[5][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n158 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[5][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[6][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n156 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[6][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[7][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n150 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[7][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[8][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n148 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[8][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[9][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n146 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[9][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[10][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n144 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[10][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[11][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n142 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[11][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[12][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n140 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[12][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[13][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n138 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[13][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[14][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n136 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[14][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[15][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n133 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[15][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[16][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n131 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[16][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[17][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n129 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[17][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[18][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n127 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[18][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[19][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n125 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[19][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[20][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n123 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[20][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[21][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n121 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[21][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[22][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n119 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[22][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[23][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n116 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[23][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[25][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n112 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[25][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[26][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n110 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[26][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[27][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n108 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[27][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[28][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n106 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[28][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[29][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n104 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[29][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[30][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n102 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[30][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[31][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n99 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[31][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[32][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n97 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[32][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[33][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n95 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[33][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[34][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n93 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[34][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[35][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[35][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[36][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n89 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[36][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[37][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n87 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[37][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[38][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n85 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[38][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[39][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n82 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[39][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[40][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n80 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[40][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[41][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n78 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[41][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[42][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n76 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[42][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[43][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[43][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[44][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[44][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[45][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[45][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[46][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[46][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[47][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[47][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[48][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[48][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[49][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[49][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[50][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[50][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[51][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[51][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[52][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[52][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[53][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[53][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[54][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[54][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[55][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[55][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[56][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[56][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[57][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[57][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[58][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[58][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[59][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[59][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[60][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[60][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[61][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[61][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[62][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[62][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[63][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[63][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[24][4]  ( .D(\i_fifo_rx/n7 ), .E(\i_fifo_rx/n114 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[24][4] ) );
  DFEC1 \i_fifo_rx/mem_reg[0][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n168 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[0][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[1][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n166 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[1][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[2][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n164 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[2][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[3][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n162 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[3][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[4][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n160 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[4][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[5][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n158 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[5][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[6][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n156 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[6][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[7][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n150 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[7][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[8][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n148 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[8][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[9][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n146 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[9][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[10][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n144 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[10][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[11][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n142 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[11][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[12][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n140 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[12][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[13][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n138 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[13][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[14][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n136 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[14][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[15][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n133 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[15][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[16][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n131 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[16][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[17][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n129 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[17][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[18][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n127 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[18][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[19][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n125 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[19][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[20][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n123 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[20][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[21][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n121 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[21][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[22][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n119 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[22][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[23][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n116 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[23][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[25][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n112 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[25][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[26][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n110 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[26][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[27][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n108 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[27][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[28][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n106 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[28][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[29][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n104 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[29][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[30][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n102 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[30][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[31][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n99 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[31][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[32][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n97 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[32][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[33][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n95 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[33][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[34][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n93 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[34][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[35][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[35][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[36][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n89 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[36][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[37][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n87 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[37][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[38][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n85 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[38][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[39][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n82 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[39][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[40][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n80 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[40][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[41][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n78 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[41][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[42][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n76 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[42][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[43][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[43][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[44][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[44][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[45][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[45][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[46][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[46][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[47][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[47][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[48][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[48][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[49][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[49][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[50][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[50][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[51][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[51][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[52][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[52][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[53][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[53][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[54][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[54][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[55][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[55][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[56][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[56][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[57][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[57][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[58][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[58][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[59][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[59][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[60][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[60][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[61][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[61][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[62][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[62][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[63][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[63][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[24][5]  ( .D(\i_fifo_rx/n8 ), .E(\i_fifo_rx/n114 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[24][5] ) );
  DFEC1 \i_fifo_rx/mem_reg[0][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n168 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[0][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[1][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n166 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[1][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[2][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n164 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[2][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[3][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n162 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[3][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[4][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n160 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[4][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[5][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n158 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[5][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[6][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n156 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[6][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[7][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n150 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[7][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[8][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n148 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[8][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[9][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n146 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[9][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[10][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n144 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[10][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[11][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n142 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[11][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[12][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n140 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[12][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[13][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n138 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[13][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[14][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n136 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[14][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[15][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n133 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[15][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[16][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n131 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[16][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[17][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n129 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[17][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[18][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n127 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[18][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[19][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n125 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[19][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[20][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n123 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[20][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[21][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n121 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[21][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[22][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n119 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[22][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[23][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n116 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[23][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[25][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n112 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[25][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[26][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n110 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[26][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[27][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n108 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[27][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[28][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n106 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[28][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[29][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n104 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[29][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[30][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n102 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[30][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[31][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n99 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[31][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[32][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n97 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[32][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[33][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n95 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[33][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[34][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n93 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[34][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[35][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[35][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[36][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n89 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[36][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[37][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n87 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[37][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[38][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n85 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[38][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[39][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n82 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[39][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[40][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n80 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[40][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[41][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n78 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[41][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[42][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n76 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[42][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[43][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[43][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[44][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[44][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[45][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[45][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[46][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[46][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[47][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[47][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[48][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[48][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[49][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[49][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[50][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[50][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[51][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[51][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[52][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[52][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[53][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[53][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[54][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[54][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[55][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[55][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[56][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[56][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[57][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[57][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[58][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[58][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[59][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[59][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[60][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[60][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[61][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[61][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[62][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[62][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[63][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[63][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[24][6]  ( .D(\i_fifo_rx/n9 ), .E(\i_fifo_rx/n114 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[24][6] ) );
  DFEC1 \i_fifo_rx/mem_reg[0][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n168 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[0][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[1][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n166 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[1][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[2][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n164 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[2][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[3][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n162 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[3][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[4][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n160 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[4][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[5][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n158 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[5][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[6][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n156 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[6][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[7][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n150 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[7][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[8][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n148 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[8][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[9][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n146 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[9][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[10][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n144 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[10][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[11][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n142 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[11][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[12][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n140 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[12][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[13][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n138 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[13][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[14][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n136 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[14][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[15][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n133 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[15][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[16][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n131 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[16][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[17][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n129 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[17][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[18][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n127 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[18][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[19][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n125 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[19][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[20][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n123 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[20][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[21][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n121 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[21][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[22][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n119 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[22][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[23][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n116 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[23][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[25][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n112 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[25][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[26][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n110 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[26][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[27][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n108 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[27][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[28][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n106 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[28][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[29][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n104 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[29][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[30][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n102 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[30][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[31][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n99 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[31][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[32][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n97 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[32][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[33][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n95 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[33][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[34][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n93 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[34][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[35][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n91 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[35][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[36][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n89 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[36][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[37][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n87 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[37][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[38][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n85 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[38][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[39][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n82 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[39][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[40][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n80 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[40][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[41][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n78 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[41][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[42][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n76 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[42][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[43][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n74 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[43][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[44][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n72 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[44][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[45][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n70 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[45][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[46][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n68 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[46][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[47][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n65 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[47][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[48][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n63 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[48][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[49][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n61 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[49][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[50][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n59 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[50][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[51][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n57 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[51][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[52][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n55 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[52][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[53][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n53 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[53][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[54][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n51 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[54][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[55][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n48 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[55][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[56][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n42 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[56][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[57][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n39 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[57][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[58][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n36 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[58][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[59][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n33 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[59][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[60][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n30 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[60][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[61][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n27 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[61][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[62][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n24 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[62][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[63][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n12 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[63][7] ) );
  DFEC1 \i_fifo_rx/mem_reg[24][7]  ( .D(\i_fifo_rx/n10 ), .E(\i_fifo_rx/n114 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/mem[24][7] ) );
  DFEC1 \i_mod_iq/fsm_mapping/cpt_old_reg[1]  ( .D(
        \i_mod_iq/fsm_mapping/cpt [1]), .E(\i_mod_iq/fsm_mapping/N259 ), .C(
        clk_i), .RN(resetn_i), .Q(\i_mod_iq/fsm_mapping/cpt_old [1]), .QN(
        \i_mod_iq/fsm_mapping/n178 ) );
  DFEC1 \i_iq_demod/gen_sin/current_state_reg[2]  ( .D(\i_iq_demod/sine_IN [1]), .E(\i_iq_demod/gen_sin/N106 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/gen_sin/current_state [2]), .QN(\i_iq_demod/gen_sin/n5 )
         );
  IMUX40 \i_fifo_rx/U228  ( .A(\i_fifo_rx/n229 ), .B(\i_fifo_rx/n230 ), .C(
        \i_fifo_rx/n231 ), .D(\i_fifo_rx/n232 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n228 ) );
  MUX41 \i_fifo_rx/U230  ( .A(\i_fifo_rx/n233 ), .B(\i_fifo_rx/n223 ), .C(
        \i_fifo_rx/n228 ), .D(\i_fifo_rx/n218 ), .S0(\i_fifo_rx/N38 ), .S1(
        \i_fifo_rx/N37 ), .Q(\i_fifo_rx/N94 ) );
  IMUX40 \i_fifo_rx/U233  ( .A(\i_fifo_rx/n249 ), .B(\i_fifo_rx/n250 ), .C(
        \i_fifo_rx/n251 ), .D(\i_fifo_rx/n252 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n248 ) );
  MUX41 \i_fifo_rx/U235  ( .A(\i_fifo_rx/n253 ), .B(\i_fifo_rx/n243 ), .C(
        \i_fifo_rx/n248 ), .D(\i_fifo_rx/n238 ), .S0(\i_fifo_rx/N38 ), .S1(
        \i_fifo_rx/N37 ), .Q(\i_fifo_rx/N93 ) );
  IMUX40 \i_fifo_rx/U238  ( .A(\i_fifo_rx/n269 ), .B(\i_fifo_rx/n270 ), .C(
        \i_fifo_rx/n271 ), .D(\i_fifo_rx/n272 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n268 ) );
  MUX41 \i_fifo_rx/U240  ( .A(\i_fifo_rx/n273 ), .B(\i_fifo_rx/n263 ), .C(
        \i_fifo_rx/n268 ), .D(\i_fifo_rx/n258 ), .S0(\i_fifo_rx/N38 ), .S1(
        \i_fifo_rx/N37 ), .Q(\i_fifo_rx/N92 ) );
  IMUX40 \i_fifo_rx/U243  ( .A(\i_fifo_rx/n289 ), .B(\i_fifo_rx/n290 ), .C(
        \i_fifo_rx/n291 ), .D(\i_fifo_rx/n292 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n288 ) );
  MUX41 \i_fifo_rx/U245  ( .A(\i_fifo_rx/n293 ), .B(\i_fifo_rx/n283 ), .C(
        \i_fifo_rx/n288 ), .D(\i_fifo_rx/n278 ), .S0(\i_fifo_rx/N38 ), .S1(
        \i_fifo_rx/N37 ), .Q(\i_fifo_rx/N91 ) );
  IMUX40 \i_fifo_rx/U248  ( .A(\i_fifo_rx/n309 ), .B(\i_fifo_rx/n310 ), .C(
        \i_fifo_rx/n311 ), .D(\i_fifo_rx/n312 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n308 ) );
  MUX41 \i_fifo_rx/U250  ( .A(\i_fifo_rx/n313 ), .B(\i_fifo_rx/n303 ), .C(
        \i_fifo_rx/n308 ), .D(\i_fifo_rx/n298 ), .S0(\i_fifo_rx/N38 ), .S1(
        \i_fifo_rx/N37 ), .Q(\i_fifo_rx/N90 ) );
  IMUX40 \i_fifo_rx/U253  ( .A(\i_fifo_rx/n329 ), .B(\i_fifo_rx/n330 ), .C(
        \i_fifo_rx/n331 ), .D(\i_fifo_rx/n332 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n328 ) );
  MUX41 \i_fifo_rx/U255  ( .A(\i_fifo_rx/n333 ), .B(\i_fifo_rx/n323 ), .C(
        \i_fifo_rx/n328 ), .D(\i_fifo_rx/n318 ), .S0(\i_fifo_rx/N38 ), .S1(
        \i_fifo_rx/N37 ), .Q(\i_fifo_rx/N89 ) );
  IMUX40 \i_fifo_rx/U258  ( .A(\i_fifo_rx/n349 ), .B(\i_fifo_rx/n350 ), .C(
        \i_fifo_rx/n351 ), .D(\i_fifo_rx/n352 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n348 ) );
  MUX41 \i_fifo_rx/U260  ( .A(\i_fifo_rx/n353 ), .B(\i_fifo_rx/n343 ), .C(
        \i_fifo_rx/n348 ), .D(\i_fifo_rx/n338 ), .S0(\i_fifo_rx/N38 ), .S1(
        \i_fifo_rx/N37 ), .Q(\i_fifo_rx/N88 ) );
  IMUX40 \i_fifo_rx/U263  ( .A(\i_fifo_rx/n369 ), .B(\i_fifo_rx/n370 ), .C(
        \i_fifo_rx/n371 ), .D(\i_fifo_rx/n372 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n368 ) );
  MUX41 \i_fifo_rx/U265  ( .A(\i_fifo_rx/n373 ), .B(\i_fifo_rx/n363 ), .C(
        \i_fifo_rx/n368 ), .D(\i_fifo_rx/n358 ), .S0(\i_fifo_rx/N38 ), .S1(
        \i_fifo_rx/N37 ), .Q(\i_fifo_rx/N87 ) );
  IMUX40 \i_fifo_tx/U255  ( .A(\i_fifo_tx/mem[24][0] ), .B(
        \i_fifo_tx/mem[25][0] ), .C(\i_fifo_tx/mem[26][0] ), .D(
        \i_fifo_tx/mem[27][0] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n220 ) );
  IMUX40 \i_fifo_tx/U257  ( .A(\i_fifo_tx/mem[16][0] ), .B(
        \i_fifo_tx/mem[17][0] ), .C(\i_fifo_tx/mem[18][0] ), .D(
        \i_fifo_tx/mem[19][0] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n219 ) );
  IMUX40 \i_fifo_tx/U256  ( .A(\i_fifo_tx/mem[20][0] ), .B(
        \i_fifo_tx/mem[21][0] ), .C(\i_fifo_tx/mem[22][0] ), .D(
        \i_fifo_tx/mem[23][0] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n221 ) );
  IMUX40 \i_fifo_tx/U208  ( .A(\i_fifo_tx/n219 ), .B(\i_fifo_tx/n220 ), .C(
        \i_fifo_tx/n221 ), .D(\i_fifo_tx/n222 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n218 ) );
  IMUX40 \i_fifo_tx/U259  ( .A(\i_fifo_tx/mem[8][0] ), .B(
        \i_fifo_tx/mem[9][0] ), .C(\i_fifo_tx/mem[10][0] ), .D(
        \i_fifo_tx/mem[11][0] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n225 ) );
  IMUX40 \i_fifo_tx/U261  ( .A(\i_fifo_tx/mem[0][0] ), .B(
        \i_fifo_tx/mem[1][0] ), .C(\i_fifo_tx/mem[2][0] ), .D(
        \i_fifo_tx/mem[3][0] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n224 ) );
  IMUX40 \i_fifo_tx/U260  ( .A(\i_fifo_tx/mem[4][0] ), .B(
        \i_fifo_tx/mem[5][0] ), .C(\i_fifo_tx/mem[6][0] ), .D(
        \i_fifo_tx/mem[7][0] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n226 ) );
  IMUX40 \i_fifo_tx/U209  ( .A(\i_fifo_tx/n224 ), .B(\i_fifo_tx/n225 ), .C(
        \i_fifo_tx/n226 ), .D(\i_fifo_tx/n227 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n223 ) );
  IMUX40 \i_fifo_tx/U251  ( .A(\i_fifo_tx/mem[40][0] ), .B(
        \i_fifo_tx/mem[41][0] ), .C(\i_fifo_tx/mem[42][0] ), .D(
        \i_fifo_tx/mem[43][0] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n215 ) );
  IMUX40 \i_fifo_tx/U253  ( .A(\i_fifo_tx/mem[32][0] ), .B(
        \i_fifo_tx/mem[33][0] ), .C(\i_fifo_tx/mem[34][0] ), .D(
        \i_fifo_tx/mem[35][0] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n214 ) );
  IMUX40 \i_fifo_tx/U252  ( .A(\i_fifo_tx/mem[36][0] ), .B(
        \i_fifo_tx/mem[37][0] ), .C(\i_fifo_tx/mem[38][0] ), .D(
        \i_fifo_tx/mem[39][0] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n216 ) );
  IMUX40 \i_fifo_tx/U207  ( .A(\i_fifo_tx/n214 ), .B(\i_fifo_tx/n215 ), .C(
        \i_fifo_tx/n216 ), .D(\i_fifo_tx/n217 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n213 ) );
  IMUX40 \i_fifo_tx/U247  ( .A(\i_fifo_tx/mem[56][0] ), .B(
        \i_fifo_tx/mem[57][0] ), .C(\i_fifo_tx/mem[58][0] ), .D(
        \i_fifo_tx/mem[59][0] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n210 ) );
  IMUX40 \i_fifo_tx/U249  ( .A(\i_fifo_tx/mem[48][0] ), .B(
        \i_fifo_tx/mem[49][0] ), .C(\i_fifo_tx/mem[50][0] ), .D(
        \i_fifo_tx/mem[51][0] ), .S0(n317), .S1(n319), .Q(\i_fifo_tx/n209 ) );
  IMUX40 \i_fifo_tx/U248  ( .A(\i_fifo_tx/mem[52][0] ), .B(
        \i_fifo_tx/mem[53][0] ), .C(\i_fifo_tx/mem[54][0] ), .D(
        \i_fifo_tx/mem[55][0] ), .S0(n317), .S1(n319), .Q(\i_fifo_tx/n211 ) );
  IMUX40 \i_fifo_tx/U206  ( .A(\i_fifo_tx/n209 ), .B(\i_fifo_tx/n210 ), .C(
        \i_fifo_tx/n211 ), .D(\i_fifo_tx/n212 ), .S0(\i_fifo_tx/N27 ), .S1(
        n1946), .Q(\i_fifo_tx/n208 ) );
  IMUX40 \i_fifo_tx/U271  ( .A(\i_fifo_tx/mem[24][1] ), .B(
        \i_fifo_tx/mem[25][1] ), .C(\i_fifo_tx/mem[26][1] ), .D(
        \i_fifo_tx/mem[27][1] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n240 ) );
  IMUX40 \i_fifo_tx/U273  ( .A(\i_fifo_tx/mem[16][1] ), .B(
        \i_fifo_tx/mem[17][1] ), .C(\i_fifo_tx/mem[18][1] ), .D(
        \i_fifo_tx/mem[19][1] ), .S0(n317), .S1(n319), .Q(\i_fifo_tx/n239 ) );
  IMUX40 \i_fifo_tx/U272  ( .A(\i_fifo_tx/mem[20][1] ), .B(
        \i_fifo_tx/mem[21][1] ), .C(\i_fifo_tx/mem[22][1] ), .D(
        \i_fifo_tx/mem[23][1] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n241 ) );
  IMUX40 \i_fifo_tx/U213  ( .A(\i_fifo_tx/n239 ), .B(\i_fifo_tx/n240 ), .C(
        \i_fifo_tx/n241 ), .D(\i_fifo_tx/n242 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n238 ) );
  IMUX40 \i_fifo_tx/U275  ( .A(\i_fifo_tx/mem[8][1] ), .B(
        \i_fifo_tx/mem[9][1] ), .C(\i_fifo_tx/mem[10][1] ), .D(
        \i_fifo_tx/mem[11][1] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n245 ) );
  IMUX40 \i_fifo_tx/U277  ( .A(\i_fifo_tx/mem[0][1] ), .B(
        \i_fifo_tx/mem[1][1] ), .C(\i_fifo_tx/mem[2][1] ), .D(
        \i_fifo_tx/mem[3][1] ), .S0(n314), .S1(n318), .Q(\i_fifo_tx/n244 ) );
  IMUX40 \i_fifo_tx/U276  ( .A(\i_fifo_tx/mem[4][1] ), .B(
        \i_fifo_tx/mem[5][1] ), .C(\i_fifo_tx/mem[6][1] ), .D(
        \i_fifo_tx/mem[7][1] ), .S0(n317), .S1(n319), .Q(\i_fifo_tx/n246 ) );
  IMUX40 \i_fifo_tx/U214  ( .A(\i_fifo_tx/n244 ), .B(\i_fifo_tx/n245 ), .C(
        \i_fifo_tx/n246 ), .D(\i_fifo_tx/n247 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n243 ) );
  IMUX40 \i_fifo_tx/U267  ( .A(\i_fifo_tx/mem[40][1] ), .B(
        \i_fifo_tx/mem[41][1] ), .C(\i_fifo_tx/mem[42][1] ), .D(
        \i_fifo_tx/mem[43][1] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n235 ) );
  IMUX40 \i_fifo_tx/U269  ( .A(\i_fifo_tx/mem[32][1] ), .B(
        \i_fifo_tx/mem[33][1] ), .C(\i_fifo_tx/mem[34][1] ), .D(
        \i_fifo_tx/mem[35][1] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n234 ) );
  IMUX40 \i_fifo_tx/U268  ( .A(\i_fifo_tx/mem[36][1] ), .B(
        \i_fifo_tx/mem[37][1] ), .C(\i_fifo_tx/mem[38][1] ), .D(
        \i_fifo_tx/mem[39][1] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n236 ) );
  IMUX40 \i_fifo_tx/U212  ( .A(\i_fifo_tx/n234 ), .B(\i_fifo_tx/n235 ), .C(
        \i_fifo_tx/n236 ), .D(\i_fifo_tx/n237 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n233 ) );
  IMUX40 \i_fifo_tx/U263  ( .A(\i_fifo_tx/mem[56][1] ), .B(
        \i_fifo_tx/mem[57][1] ), .C(\i_fifo_tx/mem[58][1] ), .D(
        \i_fifo_tx/mem[59][1] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n230 ) );
  IMUX40 \i_fifo_tx/U265  ( .A(\i_fifo_tx/mem[48][1] ), .B(
        \i_fifo_tx/mem[49][1] ), .C(\i_fifo_tx/mem[50][1] ), .D(
        \i_fifo_tx/mem[51][1] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n229 ) );
  IMUX40 \i_fifo_tx/U264  ( .A(\i_fifo_tx/mem[52][1] ), .B(
        \i_fifo_tx/mem[53][1] ), .C(\i_fifo_tx/mem[54][1] ), .D(
        \i_fifo_tx/mem[55][1] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n231 ) );
  IMUX40 \i_fifo_tx/U211  ( .A(\i_fifo_tx/n229 ), .B(\i_fifo_tx/n230 ), .C(
        \i_fifo_tx/n231 ), .D(\i_fifo_tx/n232 ), .S0(\i_fifo_tx/N27 ), .S1(
        \i_fifo_tx/N26 ), .Q(\i_fifo_tx/n228 ) );
  IMUX40 \i_fifo_tx/U287  ( .A(\i_fifo_tx/mem[24][2] ), .B(
        \i_fifo_tx/mem[25][2] ), .C(\i_fifo_tx/mem[26][2] ), .D(
        \i_fifo_tx/mem[27][2] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n260 ) );
  IMUX40 \i_fifo_tx/U289  ( .A(\i_fifo_tx/mem[16][2] ), .B(
        \i_fifo_tx/mem[17][2] ), .C(\i_fifo_tx/mem[18][2] ), .D(
        \i_fifo_tx/mem[19][2] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n259 ) );
  IMUX40 \i_fifo_tx/U288  ( .A(\i_fifo_tx/mem[20][2] ), .B(
        \i_fifo_tx/mem[21][2] ), .C(\i_fifo_tx/mem[22][2] ), .D(
        \i_fifo_tx/mem[23][2] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n261 ) );
  IMUX40 \i_fifo_tx/U218  ( .A(\i_fifo_tx/n259 ), .B(\i_fifo_tx/n260 ), .C(
        \i_fifo_tx/n261 ), .D(\i_fifo_tx/n262 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n258 ) );
  IMUX40 \i_fifo_tx/U291  ( .A(\i_fifo_tx/mem[8][2] ), .B(
        \i_fifo_tx/mem[9][2] ), .C(\i_fifo_tx/mem[10][2] ), .D(
        \i_fifo_tx/mem[11][2] ), .S0(n314), .S1(n318), .Q(\i_fifo_tx/n265 ) );
  IMUX40 \i_fifo_tx/U293  ( .A(\i_fifo_tx/mem[0][2] ), .B(
        \i_fifo_tx/mem[1][2] ), .C(\i_fifo_tx/mem[2][2] ), .D(
        \i_fifo_tx/mem[3][2] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n264 ) );
  IMUX40 \i_fifo_tx/U292  ( .A(\i_fifo_tx/mem[4][2] ), .B(
        \i_fifo_tx/mem[5][2] ), .C(\i_fifo_tx/mem[6][2] ), .D(
        \i_fifo_tx/mem[7][2] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n266 ) );
  IMUX40 \i_fifo_tx/U219  ( .A(\i_fifo_tx/n264 ), .B(\i_fifo_tx/n265 ), .C(
        \i_fifo_tx/n266 ), .D(\i_fifo_tx/n267 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n263 ) );
  IMUX40 \i_fifo_tx/U283  ( .A(\i_fifo_tx/mem[40][2] ), .B(
        \i_fifo_tx/mem[41][2] ), .C(\i_fifo_tx/mem[42][2] ), .D(
        \i_fifo_tx/mem[43][2] ), .S0(n314), .S1(n318), .Q(\i_fifo_tx/n255 ) );
  IMUX40 \i_fifo_tx/U285  ( .A(\i_fifo_tx/mem[32][2] ), .B(
        \i_fifo_tx/mem[33][2] ), .C(\i_fifo_tx/mem[34][2] ), .D(
        \i_fifo_tx/mem[35][2] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n254 ) );
  IMUX40 \i_fifo_tx/U284  ( .A(\i_fifo_tx/mem[36][2] ), .B(
        \i_fifo_tx/mem[37][2] ), .C(\i_fifo_tx/mem[38][2] ), .D(
        \i_fifo_tx/mem[39][2] ), .S0(n132), .S1(n318), .Q(\i_fifo_tx/n256 ) );
  IMUX40 \i_fifo_tx/U217  ( .A(\i_fifo_tx/n254 ), .B(\i_fifo_tx/n255 ), .C(
        \i_fifo_tx/n256 ), .D(\i_fifo_tx/n257 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n253 ) );
  IMUX40 \i_fifo_tx/U279  ( .A(\i_fifo_tx/mem[56][2] ), .B(
        \i_fifo_tx/mem[57][2] ), .C(\i_fifo_tx/mem[58][2] ), .D(
        \i_fifo_tx/mem[59][2] ), .S0(n132), .S1(n318), .Q(\i_fifo_tx/n250 ) );
  IMUX40 \i_fifo_tx/U281  ( .A(\i_fifo_tx/mem[48][2] ), .B(
        \i_fifo_tx/mem[49][2] ), .C(\i_fifo_tx/mem[50][2] ), .D(
        \i_fifo_tx/mem[51][2] ), .S0(n314), .S1(n318), .Q(\i_fifo_tx/n249 ) );
  IMUX40 \i_fifo_tx/U280  ( .A(\i_fifo_tx/mem[52][2] ), .B(
        \i_fifo_tx/mem[53][2] ), .C(\i_fifo_tx/mem[54][2] ), .D(
        \i_fifo_tx/mem[55][2] ), .S0(n132), .S1(n318), .Q(\i_fifo_tx/n251 ) );
  IMUX40 \i_fifo_tx/U216  ( .A(\i_fifo_tx/n249 ), .B(\i_fifo_tx/n250 ), .C(
        \i_fifo_tx/n251 ), .D(\i_fifo_tx/n252 ), .S0(\i_fifo_tx/N27 ), .S1(
        \i_fifo_tx/N26 ), .Q(\i_fifo_tx/n248 ) );
  IMUX40 \i_fifo_tx/U303  ( .A(\i_fifo_tx/mem[24][3] ), .B(
        \i_fifo_tx/mem[25][3] ), .C(\i_fifo_tx/mem[26][3] ), .D(
        \i_fifo_tx/mem[27][3] ), .S0(n317), .S1(n319), .Q(\i_fifo_tx/n280 ) );
  IMUX40 \i_fifo_tx/U305  ( .A(\i_fifo_tx/mem[16][3] ), .B(
        \i_fifo_tx/mem[17][3] ), .C(\i_fifo_tx/mem[18][3] ), .D(
        \i_fifo_tx/mem[19][3] ), .S0(n317), .S1(n319), .Q(\i_fifo_tx/n279 ) );
  IMUX40 \i_fifo_tx/U304  ( .A(\i_fifo_tx/mem[20][3] ), .B(
        \i_fifo_tx/mem[21][3] ), .C(\i_fifo_tx/mem[22][3] ), .D(
        \i_fifo_tx/mem[23][3] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n281 ) );
  IMUX40 \i_fifo_tx/U223  ( .A(\i_fifo_tx/n279 ), .B(\i_fifo_tx/n280 ), .C(
        \i_fifo_tx/n281 ), .D(\i_fifo_tx/n282 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n278 ) );
  IMUX40 \i_fifo_tx/U307  ( .A(\i_fifo_tx/mem[8][3] ), .B(
        \i_fifo_tx/mem[9][3] ), .C(\i_fifo_tx/mem[10][3] ), .D(
        \i_fifo_tx/mem[11][3] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n285 ) );
  IMUX40 \i_fifo_tx/U309  ( .A(\i_fifo_tx/mem[0][3] ), .B(
        \i_fifo_tx/mem[1][3] ), .C(\i_fifo_tx/mem[2][3] ), .D(
        \i_fifo_tx/mem[3][3] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n284 ) );
  IMUX40 \i_fifo_tx/U308  ( .A(\i_fifo_tx/mem[4][3] ), .B(
        \i_fifo_tx/mem[5][3] ), .C(\i_fifo_tx/mem[6][3] ), .D(
        \i_fifo_tx/mem[7][3] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n286 ) );
  IMUX40 \i_fifo_tx/U224  ( .A(\i_fifo_tx/n284 ), .B(\i_fifo_tx/n285 ), .C(
        \i_fifo_tx/n286 ), .D(\i_fifo_tx/n287 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n283 ) );
  IMUX40 \i_fifo_tx/U299  ( .A(\i_fifo_tx/mem[40][3] ), .B(
        \i_fifo_tx/mem[41][3] ), .C(\i_fifo_tx/mem[42][3] ), .D(
        \i_fifo_tx/mem[43][3] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n275 ) );
  IMUX40 \i_fifo_tx/U301  ( .A(\i_fifo_tx/mem[32][3] ), .B(
        \i_fifo_tx/mem[33][3] ), .C(\i_fifo_tx/mem[34][3] ), .D(
        \i_fifo_tx/mem[35][3] ), .S0(n317), .S1(n319), .Q(\i_fifo_tx/n274 ) );
  IMUX40 \i_fifo_tx/U300  ( .A(\i_fifo_tx/mem[36][3] ), .B(
        \i_fifo_tx/mem[37][3] ), .C(\i_fifo_tx/mem[38][3] ), .D(
        \i_fifo_tx/mem[39][3] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n276 ) );
  IMUX40 \i_fifo_tx/U222  ( .A(\i_fifo_tx/n274 ), .B(\i_fifo_tx/n275 ), .C(
        \i_fifo_tx/n276 ), .D(\i_fifo_tx/n277 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n273 ) );
  IMUX40 \i_fifo_tx/U295  ( .A(\i_fifo_tx/mem[56][3] ), .B(
        \i_fifo_tx/mem[57][3] ), .C(\i_fifo_tx/mem[58][3] ), .D(
        \i_fifo_tx/mem[59][3] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n270 ) );
  IMUX40 \i_fifo_tx/U297  ( .A(\i_fifo_tx/mem[48][3] ), .B(
        \i_fifo_tx/mem[49][3] ), .C(\i_fifo_tx/mem[50][3] ), .D(
        \i_fifo_tx/mem[51][3] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n269 ) );
  IMUX40 \i_fifo_tx/U296  ( .A(\i_fifo_tx/mem[52][3] ), .B(
        \i_fifo_tx/mem[53][3] ), .C(\i_fifo_tx/mem[54][3] ), .D(
        \i_fifo_tx/mem[55][3] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n271 ) );
  IMUX40 \i_fifo_tx/U221  ( .A(\i_fifo_tx/n269 ), .B(\i_fifo_tx/n270 ), .C(
        \i_fifo_tx/n271 ), .D(\i_fifo_tx/n272 ), .S0(\i_fifo_tx/N27 ), .S1(
        n1946), .Q(\i_fifo_tx/n268 ) );
  IMUX40 \i_fifo_tx/U319  ( .A(\i_fifo_tx/mem[24][4] ), .B(
        \i_fifo_tx/mem[25][4] ), .C(\i_fifo_tx/mem[26][4] ), .D(
        \i_fifo_tx/mem[27][4] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n300 ) );
  IMUX40 \i_fifo_tx/U321  ( .A(\i_fifo_tx/mem[16][4] ), .B(
        \i_fifo_tx/mem[17][4] ), .C(\i_fifo_tx/mem[18][4] ), .D(
        \i_fifo_tx/mem[19][4] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n299 ) );
  IMUX40 \i_fifo_tx/U320  ( .A(\i_fifo_tx/mem[20][4] ), .B(
        \i_fifo_tx/mem[21][4] ), .C(\i_fifo_tx/mem[22][4] ), .D(
        \i_fifo_tx/mem[23][4] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n301 ) );
  IMUX40 \i_fifo_tx/U228  ( .A(\i_fifo_tx/n299 ), .B(\i_fifo_tx/n300 ), .C(
        \i_fifo_tx/n301 ), .D(\i_fifo_tx/n302 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n298 ) );
  IMUX40 \i_fifo_tx/U323  ( .A(\i_fifo_tx/mem[8][4] ), .B(
        \i_fifo_tx/mem[9][4] ), .C(\i_fifo_tx/mem[10][4] ), .D(
        \i_fifo_tx/mem[11][4] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n305 ) );
  IMUX40 \i_fifo_tx/U325  ( .A(\i_fifo_tx/mem[0][4] ), .B(
        \i_fifo_tx/mem[1][4] ), .C(\i_fifo_tx/mem[2][4] ), .D(
        \i_fifo_tx/mem[3][4] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n304 ) );
  IMUX40 \i_fifo_tx/U324  ( .A(\i_fifo_tx/mem[4][4] ), .B(
        \i_fifo_tx/mem[5][4] ), .C(\i_fifo_tx/mem[6][4] ), .D(
        \i_fifo_tx/mem[7][4] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n306 ) );
  IMUX40 \i_fifo_tx/U229  ( .A(\i_fifo_tx/n304 ), .B(\i_fifo_tx/n305 ), .C(
        \i_fifo_tx/n306 ), .D(\i_fifo_tx/n307 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n303 ) );
  IMUX40 \i_fifo_tx/U315  ( .A(\i_fifo_tx/mem[40][4] ), .B(
        \i_fifo_tx/mem[41][4] ), .C(\i_fifo_tx/mem[42][4] ), .D(
        \i_fifo_tx/mem[43][4] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n295 ) );
  IMUX40 \i_fifo_tx/U317  ( .A(\i_fifo_tx/mem[32][4] ), .B(
        \i_fifo_tx/mem[33][4] ), .C(\i_fifo_tx/mem[34][4] ), .D(
        \i_fifo_tx/mem[35][4] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n294 ) );
  IMUX40 \i_fifo_tx/U316  ( .A(\i_fifo_tx/mem[36][4] ), .B(
        \i_fifo_tx/mem[37][4] ), .C(\i_fifo_tx/mem[38][4] ), .D(
        \i_fifo_tx/mem[39][4] ), .S0(n132), .S1(n318), .Q(\i_fifo_tx/n296 ) );
  IMUX40 \i_fifo_tx/U227  ( .A(\i_fifo_tx/n294 ), .B(\i_fifo_tx/n295 ), .C(
        \i_fifo_tx/n296 ), .D(\i_fifo_tx/n297 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n293 ) );
  IMUX40 \i_fifo_tx/U311  ( .A(\i_fifo_tx/mem[56][4] ), .B(
        \i_fifo_tx/mem[57][4] ), .C(\i_fifo_tx/mem[58][4] ), .D(
        \i_fifo_tx/mem[59][4] ), .S0(n314), .S1(n318), .Q(\i_fifo_tx/n290 ) );
  IMUX40 \i_fifo_tx/U313  ( .A(\i_fifo_tx/mem[48][4] ), .B(
        \i_fifo_tx/mem[49][4] ), .C(\i_fifo_tx/mem[50][4] ), .D(
        \i_fifo_tx/mem[51][4] ), .S0(n314), .S1(n318), .Q(\i_fifo_tx/n289 ) );
  IMUX40 \i_fifo_tx/U312  ( .A(\i_fifo_tx/mem[52][4] ), .B(
        \i_fifo_tx/mem[53][4] ), .C(\i_fifo_tx/mem[54][4] ), .D(
        \i_fifo_tx/mem[55][4] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n291 ) );
  IMUX40 \i_fifo_tx/U226  ( .A(\i_fifo_tx/n289 ), .B(\i_fifo_tx/n290 ), .C(
        \i_fifo_tx/n291 ), .D(\i_fifo_tx/n292 ), .S0(\i_fifo_tx/N27 ), .S1(
        n1946), .Q(\i_fifo_tx/n288 ) );
  IMUX40 \i_fifo_tx/U335  ( .A(\i_fifo_tx/mem[24][5] ), .B(
        \i_fifo_tx/mem[25][5] ), .C(\i_fifo_tx/mem[26][5] ), .D(
        \i_fifo_tx/mem[27][5] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n320 ) );
  IMUX40 \i_fifo_tx/U337  ( .A(\i_fifo_tx/mem[16][5] ), .B(
        \i_fifo_tx/mem[17][5] ), .C(\i_fifo_tx/mem[18][5] ), .D(
        \i_fifo_tx/mem[19][5] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n319 ) );
  IMUX40 \i_fifo_tx/U336  ( .A(\i_fifo_tx/mem[20][5] ), .B(
        \i_fifo_tx/mem[21][5] ), .C(\i_fifo_tx/mem[22][5] ), .D(
        \i_fifo_tx/mem[23][5] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n321 ) );
  IMUX40 \i_fifo_tx/U233  ( .A(\i_fifo_tx/n319 ), .B(\i_fifo_tx/n320 ), .C(
        \i_fifo_tx/n321 ), .D(\i_fifo_tx/n322 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n318 ) );
  IMUX40 \i_fifo_tx/U339  ( .A(\i_fifo_tx/mem[8][5] ), .B(
        \i_fifo_tx/mem[9][5] ), .C(\i_fifo_tx/mem[10][5] ), .D(
        \i_fifo_tx/mem[11][5] ), .S0(n314), .S1(n318), .Q(\i_fifo_tx/n325 ) );
  IMUX40 \i_fifo_tx/U341  ( .A(\i_fifo_tx/mem[0][5] ), .B(
        \i_fifo_tx/mem[1][5] ), .C(\i_fifo_tx/mem[2][5] ), .D(
        \i_fifo_tx/mem[3][5] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n324 ) );
  IMUX40 \i_fifo_tx/U340  ( .A(\i_fifo_tx/mem[4][5] ), .B(
        \i_fifo_tx/mem[5][5] ), .C(\i_fifo_tx/mem[6][5] ), .D(
        \i_fifo_tx/mem[7][5] ), .S0(n314), .S1(n318), .Q(\i_fifo_tx/n326 ) );
  IMUX40 \i_fifo_tx/U234  ( .A(\i_fifo_tx/n324 ), .B(\i_fifo_tx/n325 ), .C(
        \i_fifo_tx/n326 ), .D(\i_fifo_tx/n327 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n323 ) );
  IMUX40 \i_fifo_tx/U331  ( .A(\i_fifo_tx/mem[40][5] ), .B(
        \i_fifo_tx/mem[41][5] ), .C(\i_fifo_tx/mem[42][5] ), .D(
        \i_fifo_tx/mem[43][5] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n315 ) );
  IMUX40 \i_fifo_tx/U333  ( .A(\i_fifo_tx/mem[32][5] ), .B(
        \i_fifo_tx/mem[33][5] ), .C(\i_fifo_tx/mem[34][5] ), .D(
        \i_fifo_tx/mem[35][5] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n314 ) );
  IMUX40 \i_fifo_tx/U332  ( .A(\i_fifo_tx/mem[36][5] ), .B(
        \i_fifo_tx/mem[37][5] ), .C(\i_fifo_tx/mem[38][5] ), .D(
        \i_fifo_tx/mem[39][5] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n316 ) );
  IMUX40 \i_fifo_tx/U232  ( .A(\i_fifo_tx/n314 ), .B(\i_fifo_tx/n315 ), .C(
        \i_fifo_tx/n316 ), .D(\i_fifo_tx/n317 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n313 ) );
  IMUX40 \i_fifo_tx/U327  ( .A(\i_fifo_tx/mem[56][5] ), .B(
        \i_fifo_tx/mem[57][5] ), .C(\i_fifo_tx/mem[58][5] ), .D(
        \i_fifo_tx/mem[59][5] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n310 ) );
  IMUX40 \i_fifo_tx/U329  ( .A(\i_fifo_tx/mem[48][5] ), .B(
        \i_fifo_tx/mem[49][5] ), .C(\i_fifo_tx/mem[50][5] ), .D(
        \i_fifo_tx/mem[51][5] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n309 ) );
  IMUX40 \i_fifo_tx/U328  ( .A(\i_fifo_tx/mem[52][5] ), .B(
        \i_fifo_tx/mem[53][5] ), .C(\i_fifo_tx/mem[54][5] ), .D(
        \i_fifo_tx/mem[55][5] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n311 ) );
  IMUX40 \i_fifo_tx/U231  ( .A(\i_fifo_tx/n309 ), .B(\i_fifo_tx/n310 ), .C(
        \i_fifo_tx/n311 ), .D(\i_fifo_tx/n312 ), .S0(\i_fifo_tx/N27 ), .S1(
        n1946), .Q(\i_fifo_tx/n308 ) );
  IMUX40 \i_fifo_tx/U351  ( .A(\i_fifo_tx/mem[24][6] ), .B(
        \i_fifo_tx/mem[25][6] ), .C(\i_fifo_tx/mem[26][6] ), .D(
        \i_fifo_tx/mem[27][6] ), .S0(n317), .S1(n319), .Q(\i_fifo_tx/n340 ) );
  IMUX40 \i_fifo_tx/U353  ( .A(\i_fifo_tx/mem[16][6] ), .B(
        \i_fifo_tx/mem[17][6] ), .C(\i_fifo_tx/mem[18][6] ), .D(
        \i_fifo_tx/mem[19][6] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n339 ) );
  IMUX40 \i_fifo_tx/U352  ( .A(\i_fifo_tx/mem[20][6] ), .B(
        \i_fifo_tx/mem[21][6] ), .C(\i_fifo_tx/mem[22][6] ), .D(
        \i_fifo_tx/mem[23][6] ), .S0(n314), .S1(n318), .Q(\i_fifo_tx/n341 ) );
  IMUX40 \i_fifo_tx/U238  ( .A(\i_fifo_tx/n339 ), .B(\i_fifo_tx/n340 ), .C(
        \i_fifo_tx/n341 ), .D(\i_fifo_tx/n342 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n338 ) );
  IMUX40 \i_fifo_tx/U355  ( .A(\i_fifo_tx/mem[8][6] ), .B(
        \i_fifo_tx/mem[9][6] ), .C(\i_fifo_tx/mem[10][6] ), .D(
        \i_fifo_tx/mem[11][6] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n345 ) );
  IMUX40 \i_fifo_tx/U357  ( .A(\i_fifo_tx/mem[0][6] ), .B(
        \i_fifo_tx/mem[1][6] ), .C(\i_fifo_tx/mem[2][6] ), .D(
        \i_fifo_tx/mem[3][6] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n344 ) );
  IMUX40 \i_fifo_tx/U356  ( .A(\i_fifo_tx/mem[4][6] ), .B(
        \i_fifo_tx/mem[5][6] ), .C(\i_fifo_tx/mem[6][6] ), .D(
        \i_fifo_tx/mem[7][6] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n346 ) );
  IMUX40 \i_fifo_tx/U239  ( .A(\i_fifo_tx/n344 ), .B(\i_fifo_tx/n345 ), .C(
        \i_fifo_tx/n346 ), .D(\i_fifo_tx/n347 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n343 ) );
  IMUX40 \i_fifo_tx/U347  ( .A(\i_fifo_tx/mem[40][6] ), .B(
        \i_fifo_tx/mem[41][6] ), .C(\i_fifo_tx/mem[42][6] ), .D(
        \i_fifo_tx/mem[43][6] ), .S0(n314), .S1(n318), .Q(\i_fifo_tx/n335 ) );
  IMUX40 \i_fifo_tx/U348  ( .A(\i_fifo_tx/mem[36][6] ), .B(
        \i_fifo_tx/mem[37][6] ), .C(\i_fifo_tx/mem[38][6] ), .D(
        \i_fifo_tx/mem[39][6] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n336 ) );
  IMUX40 \i_fifo_tx/U349  ( .A(\i_fifo_tx/mem[32][6] ), .B(
        \i_fifo_tx/mem[33][6] ), .C(\i_fifo_tx/mem[34][6] ), .D(
        \i_fifo_tx/mem[35][6] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n334 ) );
  IMUX40 \i_fifo_tx/U237  ( .A(\i_fifo_tx/n334 ), .B(\i_fifo_tx/n335 ), .C(
        \i_fifo_tx/n336 ), .D(\i_fifo_tx/n337 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n333 ) );
  IMUX40 \i_fifo_tx/U343  ( .A(\i_fifo_tx/mem[56][6] ), .B(
        \i_fifo_tx/mem[57][6] ), .C(\i_fifo_tx/mem[58][6] ), .D(
        \i_fifo_tx/mem[59][6] ), .S0(n314), .S1(n318), .Q(\i_fifo_tx/n330 ) );
  IMUX40 \i_fifo_tx/U345  ( .A(\i_fifo_tx/mem[48][6] ), .B(
        \i_fifo_tx/mem[49][6] ), .C(\i_fifo_tx/mem[50][6] ), .D(
        \i_fifo_tx/mem[51][6] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n329 ) );
  IMUX40 \i_fifo_tx/U344  ( .A(\i_fifo_tx/mem[52][6] ), .B(
        \i_fifo_tx/mem[53][6] ), .C(\i_fifo_tx/mem[54][6] ), .D(
        \i_fifo_tx/mem[55][6] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n331 ) );
  IMUX40 \i_fifo_tx/U236  ( .A(\i_fifo_tx/n329 ), .B(\i_fifo_tx/n330 ), .C(
        \i_fifo_tx/n331 ), .D(\i_fifo_tx/n332 ), .S0(\i_fifo_tx/N27 ), .S1(
        \i_fifo_tx/N26 ), .Q(\i_fifo_tx/n328 ) );
  IMUX40 \i_fifo_tx/U367  ( .A(\i_fifo_tx/mem[24][7] ), .B(
        \i_fifo_tx/mem[25][7] ), .C(\i_fifo_tx/mem[26][7] ), .D(
        \i_fifo_tx/mem[27][7] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n360 ) );
  IMUX40 \i_fifo_tx/U369  ( .A(\i_fifo_tx/mem[16][7] ), .B(
        \i_fifo_tx/mem[17][7] ), .C(\i_fifo_tx/mem[18][7] ), .D(
        \i_fifo_tx/mem[19][7] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n359 ) );
  IMUX40 \i_fifo_tx/U368  ( .A(\i_fifo_tx/mem[20][7] ), .B(
        \i_fifo_tx/mem[21][7] ), .C(\i_fifo_tx/mem[22][7] ), .D(
        \i_fifo_tx/mem[23][7] ), .S0(n317), .S1(n319), .Q(\i_fifo_tx/n361 ) );
  IMUX40 \i_fifo_tx/U243  ( .A(\i_fifo_tx/n359 ), .B(\i_fifo_tx/n360 ), .C(
        \i_fifo_tx/n361 ), .D(\i_fifo_tx/n362 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n358 ) );
  IMUX40 \i_fifo_tx/U370  ( .A(\i_fifo_tx/mem[12][7] ), .B(
        \i_fifo_tx/mem[13][7] ), .C(\i_fifo_tx/mem[14][7] ), .D(
        \i_fifo_tx/mem[15][7] ), .S0(n132), .S1(n318), .Q(\i_fifo_tx/n367 ) );
  IMUX40 \i_fifo_tx/U371  ( .A(\i_fifo_tx/mem[8][7] ), .B(
        \i_fifo_tx/mem[9][7] ), .C(\i_fifo_tx/mem[10][7] ), .D(
        \i_fifo_tx/mem[11][7] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n365 ) );
  IMUX40 \i_fifo_tx/U372  ( .A(\i_fifo_tx/mem[4][7] ), .B(
        \i_fifo_tx/mem[5][7] ), .C(\i_fifo_tx/mem[6][7] ), .D(
        \i_fifo_tx/mem[7][7] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n366 ) );
  IMUX40 \i_fifo_tx/U244  ( .A(\i_fifo_tx/n364 ), .B(\i_fifo_tx/n365 ), .C(
        \i_fifo_tx/n366 ), .D(\i_fifo_tx/n367 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n363 ) );
  IMUX40 \i_fifo_tx/U363  ( .A(\i_fifo_tx/mem[40][7] ), .B(
        \i_fifo_tx/mem[41][7] ), .C(\i_fifo_tx/mem[42][7] ), .D(
        \i_fifo_tx/mem[43][7] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n355 ) );
  IMUX40 \i_fifo_tx/U365  ( .A(\i_fifo_tx/mem[32][7] ), .B(
        \i_fifo_tx/mem[33][7] ), .C(\i_fifo_tx/mem[34][7] ), .D(
        \i_fifo_tx/mem[35][7] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n354 ) );
  IMUX40 \i_fifo_tx/U364  ( .A(\i_fifo_tx/mem[36][7] ), .B(
        \i_fifo_tx/mem[37][7] ), .C(\i_fifo_tx/mem[38][7] ), .D(
        \i_fifo_tx/mem[39][7] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n356 ) );
  IMUX40 \i_fifo_tx/U242  ( .A(\i_fifo_tx/n354 ), .B(\i_fifo_tx/n355 ), .C(
        \i_fifo_tx/n356 ), .D(\i_fifo_tx/n357 ), .S0(n273), .S1(n1946), .Q(
        \i_fifo_tx/n353 ) );
  IMUX40 \i_fifo_tx/U359  ( .A(\i_fifo_tx/mem[56][7] ), .B(
        \i_fifo_tx/mem[57][7] ), .C(\i_fifo_tx/mem[58][7] ), .D(
        \i_fifo_tx/mem[59][7] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n350 ) );
  IMUX40 \i_fifo_tx/U361  ( .A(\i_fifo_tx/mem[48][7] ), .B(
        \i_fifo_tx/mem[49][7] ), .C(\i_fifo_tx/mem[50][7] ), .D(
        \i_fifo_tx/mem[51][7] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n349 ) );
  IMUX40 \i_fifo_tx/U360  ( .A(\i_fifo_tx/mem[52][7] ), .B(
        \i_fifo_tx/mem[53][7] ), .C(\i_fifo_tx/mem[54][7] ), .D(
        \i_fifo_tx/mem[55][7] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n351 ) );
  IMUX40 \i_fifo_tx/U241  ( .A(\i_fifo_tx/n349 ), .B(\i_fifo_tx/n350 ), .C(
        \i_fifo_tx/n351 ), .D(\i_fifo_tx/n352 ), .S0(\i_fifo_tx/N27 ), .S1(
        \i_fifo_tx/N26 ), .Q(\i_fifo_tx/n348 ) );
  IMUX40 \i_fifo_rx/U447  ( .A(\i_fifo_rx/mem[8][0] ), .B(
        \i_fifo_rx/mem[9][0] ), .C(\i_fifo_rx/mem[10][0] ), .D(
        \i_fifo_rx/mem[11][0] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n395 ) );
  IMUX40 \i_fifo_rx/U449  ( .A(\i_fifo_rx/mem[0][0] ), .B(
        \i_fifo_rx/mem[1][0] ), .C(\i_fifo_rx/mem[2][0] ), .D(
        \i_fifo_rx/mem[3][0] ), .S0(n307), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n394 ) );
  IMUX40 \i_fifo_rx/U448  ( .A(\i_fifo_rx/mem[4][0] ), .B(
        \i_fifo_rx/mem[5][0] ), .C(\i_fifo_rx/mem[6][0] ), .D(
        \i_fifo_rx/mem[7][0] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n396 ) );
  IMUX40 \i_fifo_rx/U397  ( .A(\i_fifo_rx/n394 ), .B(\i_fifo_rx/n395 ), .C(
        \i_fifo_rx/n396 ), .D(\i_fifo_rx/n397 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n393 ) );
  IMUX40 \i_fifo_rx/U439  ( .A(\i_fifo_rx/mem[40][0] ), .B(
        \i_fifo_rx/mem[41][0] ), .C(\i_fifo_rx/mem[42][0] ), .D(
        \i_fifo_rx/mem[43][0] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n385 ) );
  IMUX40 \i_fifo_rx/U441  ( .A(\i_fifo_rx/mem[32][0] ), .B(
        \i_fifo_rx/mem[33][0] ), .C(\i_fifo_rx/mem[34][0] ), .D(
        \i_fifo_rx/mem[35][0] ), .S0(n307), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n384 ) );
  IMUX40 \i_fifo_rx/U440  ( .A(\i_fifo_rx/mem[36][0] ), .B(
        \i_fifo_rx/mem[37][0] ), .C(\i_fifo_rx/mem[38][0] ), .D(
        \i_fifo_rx/mem[39][0] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n386 ) );
  IMUX40 \i_fifo_rx/U395  ( .A(\i_fifo_rx/n384 ), .B(\i_fifo_rx/n385 ), .C(
        \i_fifo_rx/n386 ), .D(\i_fifo_rx/n387 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n383 ) );
  IMUX40 \i_fifo_rx/U435  ( .A(\i_fifo_rx/mem[56][0] ), .B(
        \i_fifo_rx/mem[57][0] ), .C(\i_fifo_rx/mem[58][0] ), .D(
        \i_fifo_rx/mem[59][0] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n380 ) );
  IMUX40 \i_fifo_rx/U437  ( .A(\i_fifo_rx/mem[48][0] ), .B(
        \i_fifo_rx/mem[49][0] ), .C(\i_fifo_rx/mem[50][0] ), .D(
        \i_fifo_rx/mem[51][0] ), .S0(n307), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n379 ) );
  IMUX40 \i_fifo_rx/U436  ( .A(\i_fifo_rx/mem[52][0] ), .B(
        \i_fifo_rx/mem[53][0] ), .C(\i_fifo_rx/mem[54][0] ), .D(
        \i_fifo_rx/mem[55][0] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n381 ) );
  IMUX40 \i_fifo_rx/U394  ( .A(\i_fifo_rx/n379 ), .B(\i_fifo_rx/n380 ), .C(
        \i_fifo_rx/n381 ), .D(\i_fifo_rx/n382 ), .S0(\i_fifo_rx/N42 ), .S1(
        n1939), .Q(\i_fifo_rx/n378 ) );
  IMUX40 \i_fifo_rx/U444  ( .A(\i_fifo_rx/mem[20][0] ), .B(
        \i_fifo_rx/mem[21][0] ), .C(\i_fifo_rx/mem[22][0] ), .D(
        \i_fifo_rx/mem[23][0] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n391 ) );
  IMUX40 \i_fifo_rx/U445  ( .A(\i_fifo_rx/mem[16][0] ), .B(
        \i_fifo_rx/mem[17][0] ), .C(\i_fifo_rx/mem[18][0] ), .D(
        \i_fifo_rx/mem[19][0] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n389 ) );
  IMUX40 \i_fifo_rx/U443  ( .A(\i_fifo_rx/mem[24][0] ), .B(
        \i_fifo_rx/mem[25][0] ), .C(\i_fifo_rx/mem[26][0] ), .D(
        \i_fifo_rx/mem[27][0] ), .S0(n307), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n390 ) );
  IMUX40 \i_fifo_rx/U442  ( .A(\i_fifo_rx/mem[28][0] ), .B(
        \i_fifo_rx/mem[29][0] ), .C(\i_fifo_rx/mem[30][0] ), .D(
        \i_fifo_rx/mem[31][0] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n392 ) );
  IMUX40 \i_fifo_rx/U463  ( .A(\i_fifo_rx/mem[8][1] ), .B(
        \i_fifo_rx/mem[9][1] ), .C(\i_fifo_rx/mem[10][1] ), .D(
        \i_fifo_rx/mem[11][1] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n415 ) );
  IMUX40 \i_fifo_rx/U465  ( .A(\i_fifo_rx/mem[0][1] ), .B(
        \i_fifo_rx/mem[1][1] ), .C(\i_fifo_rx/mem[2][1] ), .D(
        \i_fifo_rx/mem[3][1] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n414 ) );
  IMUX40 \i_fifo_rx/U464  ( .A(\i_fifo_rx/mem[4][1] ), .B(
        \i_fifo_rx/mem[5][1] ), .C(\i_fifo_rx/mem[6][1] ), .D(
        \i_fifo_rx/mem[7][1] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n416 ) );
  IMUX40 \i_fifo_rx/U402  ( .A(\i_fifo_rx/n414 ), .B(\i_fifo_rx/n415 ), .C(
        \i_fifo_rx/n416 ), .D(\i_fifo_rx/n417 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n413 ) );
  IMUX40 \i_fifo_rx/U455  ( .A(\i_fifo_rx/mem[40][1] ), .B(
        \i_fifo_rx/mem[41][1] ), .C(\i_fifo_rx/mem[42][1] ), .D(
        \i_fifo_rx/mem[43][1] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n405 ) );
  IMUX40 \i_fifo_rx/U457  ( .A(\i_fifo_rx/mem[32][1] ), .B(
        \i_fifo_rx/mem[33][1] ), .C(\i_fifo_rx/mem[34][1] ), .D(
        \i_fifo_rx/mem[35][1] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n404 ) );
  IMUX40 \i_fifo_rx/U456  ( .A(\i_fifo_rx/mem[36][1] ), .B(
        \i_fifo_rx/mem[37][1] ), .C(\i_fifo_rx/mem[38][1] ), .D(
        \i_fifo_rx/mem[39][1] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n406 ) );
  IMUX40 \i_fifo_rx/U400  ( .A(\i_fifo_rx/n404 ), .B(\i_fifo_rx/n405 ), .C(
        \i_fifo_rx/n406 ), .D(\i_fifo_rx/n407 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n403 ) );
  IMUX40 \i_fifo_rx/U451  ( .A(\i_fifo_rx/mem[56][1] ), .B(
        \i_fifo_rx/mem[57][1] ), .C(\i_fifo_rx/mem[58][1] ), .D(
        \i_fifo_rx/mem[59][1] ), .S0(n307), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n400 ) );
  IMUX40 \i_fifo_rx/U453  ( .A(\i_fifo_rx/mem[48][1] ), .B(
        \i_fifo_rx/mem[49][1] ), .C(\i_fifo_rx/mem[50][1] ), .D(
        \i_fifo_rx/mem[51][1] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n399 ) );
  IMUX40 \i_fifo_rx/U452  ( .A(\i_fifo_rx/mem[52][1] ), .B(
        \i_fifo_rx/mem[53][1] ), .C(\i_fifo_rx/mem[54][1] ), .D(
        \i_fifo_rx/mem[55][1] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n401 ) );
  IMUX40 \i_fifo_rx/U399  ( .A(\i_fifo_rx/n399 ), .B(\i_fifo_rx/n400 ), .C(
        \i_fifo_rx/n401 ), .D(\i_fifo_rx/n402 ), .S0(\i_fifo_rx/N42 ), .S1(
        \i_fifo_rx/N41 ), .Q(\i_fifo_rx/n398 ) );
  IMUX40 \i_fifo_rx/U460  ( .A(\i_fifo_rx/mem[20][1] ), .B(
        \i_fifo_rx/mem[21][1] ), .C(\i_fifo_rx/mem[22][1] ), .D(
        \i_fifo_rx/mem[23][1] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n411 ) );
  IMUX40 \i_fifo_rx/U461  ( .A(\i_fifo_rx/mem[16][1] ), .B(
        \i_fifo_rx/mem[17][1] ), .C(\i_fifo_rx/mem[18][1] ), .D(
        \i_fifo_rx/mem[19][1] ), .S0(\i_fifo_rx/N39 ), .S1(\i_fifo_rx/N40 ), 
        .Q(\i_fifo_rx/n409 ) );
  IMUX40 \i_fifo_rx/U459  ( .A(\i_fifo_rx/mem[24][1] ), .B(
        \i_fifo_rx/mem[25][1] ), .C(\i_fifo_rx/mem[26][1] ), .D(
        \i_fifo_rx/mem[27][1] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n410 ) );
  IMUX40 \i_fifo_rx/U458  ( .A(\i_fifo_rx/mem[28][1] ), .B(
        \i_fifo_rx/mem[29][1] ), .C(\i_fifo_rx/mem[30][1] ), .D(
        \i_fifo_rx/mem[31][1] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n412 ) );
  IMUX40 \i_fifo_rx/U479  ( .A(\i_fifo_rx/mem[8][2] ), .B(
        \i_fifo_rx/mem[9][2] ), .C(\i_fifo_rx/mem[10][2] ), .D(
        \i_fifo_rx/mem[11][2] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n435 ) );
  IMUX40 \i_fifo_rx/U481  ( .A(\i_fifo_rx/mem[0][2] ), .B(
        \i_fifo_rx/mem[1][2] ), .C(\i_fifo_rx/mem[2][2] ), .D(
        \i_fifo_rx/mem[3][2] ), .S0(n307), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n434 ) );
  IMUX40 \i_fifo_rx/U480  ( .A(\i_fifo_rx/mem[4][2] ), .B(
        \i_fifo_rx/mem[5][2] ), .C(\i_fifo_rx/mem[6][2] ), .D(
        \i_fifo_rx/mem[7][2] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n436 ) );
  IMUX40 \i_fifo_rx/U407  ( .A(\i_fifo_rx/n434 ), .B(\i_fifo_rx/n435 ), .C(
        \i_fifo_rx/n436 ), .D(\i_fifo_rx/n437 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n433 ) );
  IMUX40 \i_fifo_rx/U471  ( .A(\i_fifo_rx/mem[40][2] ), .B(
        \i_fifo_rx/mem[41][2] ), .C(\i_fifo_rx/mem[42][2] ), .D(
        \i_fifo_rx/mem[43][2] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n425 ) );
  IMUX40 \i_fifo_rx/U473  ( .A(\i_fifo_rx/mem[32][2] ), .B(
        \i_fifo_rx/mem[33][2] ), .C(\i_fifo_rx/mem[34][2] ), .D(
        \i_fifo_rx/mem[35][2] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n424 ) );
  IMUX40 \i_fifo_rx/U472  ( .A(\i_fifo_rx/mem[36][2] ), .B(
        \i_fifo_rx/mem[37][2] ), .C(\i_fifo_rx/mem[38][2] ), .D(
        \i_fifo_rx/mem[39][2] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n426 ) );
  IMUX40 \i_fifo_rx/U405  ( .A(\i_fifo_rx/n424 ), .B(\i_fifo_rx/n425 ), .C(
        \i_fifo_rx/n426 ), .D(\i_fifo_rx/n427 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n423 ) );
  IMUX40 \i_fifo_rx/U467  ( .A(\i_fifo_rx/mem[56][2] ), .B(
        \i_fifo_rx/mem[57][2] ), .C(\i_fifo_rx/mem[58][2] ), .D(
        \i_fifo_rx/mem[59][2] ), .S0(\i_fifo_rx/N39 ), .S1(n311), .Q(
        \i_fifo_rx/n420 ) );
  IMUX40 \i_fifo_rx/U469  ( .A(\i_fifo_rx/mem[48][2] ), .B(
        \i_fifo_rx/mem[49][2] ), .C(\i_fifo_rx/mem[50][2] ), .D(
        \i_fifo_rx/mem[51][2] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n419 ) );
  IMUX40 \i_fifo_rx/U468  ( .A(\i_fifo_rx/mem[52][2] ), .B(
        \i_fifo_rx/mem[53][2] ), .C(\i_fifo_rx/mem[54][2] ), .D(
        \i_fifo_rx/mem[55][2] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n421 ) );
  IMUX40 \i_fifo_rx/U404  ( .A(\i_fifo_rx/n419 ), .B(\i_fifo_rx/n420 ), .C(
        \i_fifo_rx/n421 ), .D(\i_fifo_rx/n422 ), .S0(\i_fifo_rx/N42 ), .S1(
        \i_fifo_rx/N41 ), .Q(\i_fifo_rx/n418 ) );
  IMUX40 \i_fifo_rx/U476  ( .A(\i_fifo_rx/mem[20][2] ), .B(
        \i_fifo_rx/mem[21][2] ), .C(\i_fifo_rx/mem[22][2] ), .D(
        \i_fifo_rx/mem[23][2] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n431 ) );
  IMUX40 \i_fifo_rx/U477  ( .A(\i_fifo_rx/mem[16][2] ), .B(
        \i_fifo_rx/mem[17][2] ), .C(\i_fifo_rx/mem[18][2] ), .D(
        \i_fifo_rx/mem[19][2] ), .S0(n307), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n429 ) );
  IMUX40 \i_fifo_rx/U475  ( .A(\i_fifo_rx/mem[24][2] ), .B(
        \i_fifo_rx/mem[25][2] ), .C(\i_fifo_rx/mem[26][2] ), .D(
        \i_fifo_rx/mem[27][2] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n430 ) );
  IMUX40 \i_fifo_rx/U474  ( .A(\i_fifo_rx/mem[28][2] ), .B(
        \i_fifo_rx/mem[29][2] ), .C(\i_fifo_rx/mem[30][2] ), .D(
        \i_fifo_rx/mem[31][2] ), .S0(n307), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n432 ) );
  IMUX40 \i_fifo_rx/U495  ( .A(\i_fifo_rx/mem[8][3] ), .B(
        \i_fifo_rx/mem[9][3] ), .C(\i_fifo_rx/mem[10][3] ), .D(
        \i_fifo_rx/mem[11][3] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n455 ) );
  IMUX40 \i_fifo_rx/U497  ( .A(\i_fifo_rx/mem[0][3] ), .B(
        \i_fifo_rx/mem[1][3] ), .C(\i_fifo_rx/mem[2][3] ), .D(
        \i_fifo_rx/mem[3][3] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n454 ) );
  IMUX40 \i_fifo_rx/U496  ( .A(\i_fifo_rx/mem[4][3] ), .B(
        \i_fifo_rx/mem[5][3] ), .C(\i_fifo_rx/mem[6][3] ), .D(
        \i_fifo_rx/mem[7][3] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n456 ) );
  IMUX40 \i_fifo_rx/U412  ( .A(\i_fifo_rx/n454 ), .B(\i_fifo_rx/n455 ), .C(
        \i_fifo_rx/n456 ), .D(\i_fifo_rx/n457 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n453 ) );
  IMUX40 \i_fifo_rx/U487  ( .A(\i_fifo_rx/mem[40][3] ), .B(
        \i_fifo_rx/mem[41][3] ), .C(\i_fifo_rx/mem[42][3] ), .D(
        \i_fifo_rx/mem[43][3] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n445 ) );
  IMUX40 \i_fifo_rx/U489  ( .A(\i_fifo_rx/mem[32][3] ), .B(
        \i_fifo_rx/mem[33][3] ), .C(\i_fifo_rx/mem[34][3] ), .D(
        \i_fifo_rx/mem[35][3] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n444 ) );
  IMUX40 \i_fifo_rx/U488  ( .A(\i_fifo_rx/mem[36][3] ), .B(
        \i_fifo_rx/mem[37][3] ), .C(\i_fifo_rx/mem[38][3] ), .D(
        \i_fifo_rx/mem[39][3] ), .S0(n307), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n446 ) );
  IMUX40 \i_fifo_rx/U410  ( .A(\i_fifo_rx/n444 ), .B(\i_fifo_rx/n445 ), .C(
        \i_fifo_rx/n446 ), .D(\i_fifo_rx/n447 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n443 ) );
  IMUX40 \i_fifo_rx/U483  ( .A(\i_fifo_rx/mem[56][3] ), .B(
        \i_fifo_rx/mem[57][3] ), .C(\i_fifo_rx/mem[58][3] ), .D(
        \i_fifo_rx/mem[59][3] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n440 ) );
  IMUX40 \i_fifo_rx/U485  ( .A(\i_fifo_rx/mem[48][3] ), .B(
        \i_fifo_rx/mem[49][3] ), .C(\i_fifo_rx/mem[50][3] ), .D(
        \i_fifo_rx/mem[51][3] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n439 ) );
  IMUX40 \i_fifo_rx/U484  ( .A(\i_fifo_rx/mem[52][3] ), .B(
        \i_fifo_rx/mem[53][3] ), .C(\i_fifo_rx/mem[54][3] ), .D(
        \i_fifo_rx/mem[55][3] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n441 ) );
  IMUX40 \i_fifo_rx/U409  ( .A(\i_fifo_rx/n439 ), .B(\i_fifo_rx/n440 ), .C(
        \i_fifo_rx/n441 ), .D(\i_fifo_rx/n442 ), .S0(\i_fifo_rx/N42 ), .S1(
        \i_fifo_rx/N41 ), .Q(\i_fifo_rx/n438 ) );
  IMUX40 \i_fifo_rx/U492  ( .A(\i_fifo_rx/mem[20][3] ), .B(
        \i_fifo_rx/mem[21][3] ), .C(\i_fifo_rx/mem[22][3] ), .D(
        \i_fifo_rx/mem[23][3] ), .S0(n307), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n451 ) );
  IMUX40 \i_fifo_rx/U493  ( .A(\i_fifo_rx/mem[16][3] ), .B(
        \i_fifo_rx/mem[17][3] ), .C(\i_fifo_rx/mem[18][3] ), .D(
        \i_fifo_rx/mem[19][3] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n449 ) );
  IMUX40 \i_fifo_rx/U491  ( .A(\i_fifo_rx/mem[24][3] ), .B(
        \i_fifo_rx/mem[25][3] ), .C(\i_fifo_rx/mem[26][3] ), .D(
        \i_fifo_rx/mem[27][3] ), .S0(\i_fifo_rx/N39 ), .S1(n311), .Q(
        \i_fifo_rx/n450 ) );
  IMUX40 \i_fifo_rx/U490  ( .A(\i_fifo_rx/mem[28][3] ), .B(
        \i_fifo_rx/mem[29][3] ), .C(\i_fifo_rx/mem[30][3] ), .D(
        \i_fifo_rx/mem[31][3] ), .S0(n307), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n452 ) );
  IMUX40 \i_fifo_rx/U511  ( .A(\i_fifo_rx/mem[8][4] ), .B(
        \i_fifo_rx/mem[9][4] ), .C(\i_fifo_rx/mem[10][4] ), .D(
        \i_fifo_rx/mem[11][4] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n475 ) );
  IMUX40 \i_fifo_rx/U513  ( .A(\i_fifo_rx/mem[0][4] ), .B(
        \i_fifo_rx/mem[1][4] ), .C(\i_fifo_rx/mem[2][4] ), .D(
        \i_fifo_rx/mem[3][4] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n474 ) );
  IMUX40 \i_fifo_rx/U512  ( .A(\i_fifo_rx/mem[4][4] ), .B(
        \i_fifo_rx/mem[5][4] ), .C(\i_fifo_rx/mem[6][4] ), .D(
        \i_fifo_rx/mem[7][4] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n476 ) );
  IMUX40 \i_fifo_rx/U417  ( .A(\i_fifo_rx/n474 ), .B(\i_fifo_rx/n475 ), .C(
        \i_fifo_rx/n476 ), .D(\i_fifo_rx/n477 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n473 ) );
  IMUX40 \i_fifo_rx/U503  ( .A(\i_fifo_rx/mem[40][4] ), .B(
        \i_fifo_rx/mem[41][4] ), .C(\i_fifo_rx/mem[42][4] ), .D(
        \i_fifo_rx/mem[43][4] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n465 ) );
  IMUX40 \i_fifo_rx/U505  ( .A(\i_fifo_rx/mem[32][4] ), .B(
        \i_fifo_rx/mem[33][4] ), .C(\i_fifo_rx/mem[34][4] ), .D(
        \i_fifo_rx/mem[35][4] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n464 ) );
  IMUX40 \i_fifo_rx/U504  ( .A(\i_fifo_rx/mem[36][4] ), .B(
        \i_fifo_rx/mem[37][4] ), .C(\i_fifo_rx/mem[38][4] ), .D(
        \i_fifo_rx/mem[39][4] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n466 ) );
  IMUX40 \i_fifo_rx/U415  ( .A(\i_fifo_rx/n464 ), .B(\i_fifo_rx/n465 ), .C(
        \i_fifo_rx/n466 ), .D(\i_fifo_rx/n467 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n463 ) );
  IMUX40 \i_fifo_rx/U499  ( .A(\i_fifo_rx/mem[56][4] ), .B(
        \i_fifo_rx/mem[57][4] ), .C(\i_fifo_rx/mem[58][4] ), .D(
        \i_fifo_rx/mem[59][4] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n460 ) );
  IMUX40 \i_fifo_rx/U501  ( .A(\i_fifo_rx/mem[48][4] ), .B(
        \i_fifo_rx/mem[49][4] ), .C(\i_fifo_rx/mem[50][4] ), .D(
        \i_fifo_rx/mem[51][4] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n459 ) );
  IMUX40 \i_fifo_rx/U500  ( .A(\i_fifo_rx/mem[52][4] ), .B(
        \i_fifo_rx/mem[53][4] ), .C(\i_fifo_rx/mem[54][4] ), .D(
        \i_fifo_rx/mem[55][4] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n461 ) );
  IMUX40 \i_fifo_rx/U414  ( .A(\i_fifo_rx/n459 ), .B(\i_fifo_rx/n460 ), .C(
        \i_fifo_rx/n461 ), .D(\i_fifo_rx/n462 ), .S0(\i_fifo_rx/N42 ), .S1(
        \i_fifo_rx/N41 ), .Q(\i_fifo_rx/n458 ) );
  IMUX40 \i_fifo_rx/U508  ( .A(\i_fifo_rx/mem[20][4] ), .B(
        \i_fifo_rx/mem[21][4] ), .C(\i_fifo_rx/mem[22][4] ), .D(
        \i_fifo_rx/mem[23][4] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n471 ) );
  IMUX40 \i_fifo_rx/U509  ( .A(\i_fifo_rx/mem[16][4] ), .B(
        \i_fifo_rx/mem[17][4] ), .C(\i_fifo_rx/mem[18][4] ), .D(
        \i_fifo_rx/mem[19][4] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n469 ) );
  IMUX40 \i_fifo_rx/U507  ( .A(\i_fifo_rx/mem[24][4] ), .B(
        \i_fifo_rx/mem[25][4] ), .C(\i_fifo_rx/mem[26][4] ), .D(
        \i_fifo_rx/mem[27][4] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n470 ) );
  IMUX40 \i_fifo_rx/U506  ( .A(\i_fifo_rx/mem[28][4] ), .B(
        \i_fifo_rx/mem[29][4] ), .C(\i_fifo_rx/mem[30][4] ), .D(
        \i_fifo_rx/mem[31][4] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n472 ) );
  IMUX40 \i_fifo_rx/U527  ( .A(\i_fifo_rx/mem[8][5] ), .B(
        \i_fifo_rx/mem[9][5] ), .C(\i_fifo_rx/mem[10][5] ), .D(
        \i_fifo_rx/mem[11][5] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n495 ) );
  IMUX40 \i_fifo_rx/U529  ( .A(\i_fifo_rx/mem[0][5] ), .B(
        \i_fifo_rx/mem[1][5] ), .C(\i_fifo_rx/mem[2][5] ), .D(
        \i_fifo_rx/mem[3][5] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n494 ) );
  IMUX40 \i_fifo_rx/U528  ( .A(\i_fifo_rx/mem[4][5] ), .B(
        \i_fifo_rx/mem[5][5] ), .C(\i_fifo_rx/mem[6][5] ), .D(
        \i_fifo_rx/mem[7][5] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n496 ) );
  IMUX40 \i_fifo_rx/U422  ( .A(\i_fifo_rx/n494 ), .B(\i_fifo_rx/n495 ), .C(
        \i_fifo_rx/n496 ), .D(\i_fifo_rx/n497 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n493 ) );
  IMUX40 \i_fifo_rx/U519  ( .A(\i_fifo_rx/mem[40][5] ), .B(
        \i_fifo_rx/mem[41][5] ), .C(\i_fifo_rx/mem[42][5] ), .D(
        \i_fifo_rx/mem[43][5] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n485 ) );
  IMUX40 \i_fifo_rx/U521  ( .A(\i_fifo_rx/mem[32][5] ), .B(
        \i_fifo_rx/mem[33][5] ), .C(\i_fifo_rx/mem[34][5] ), .D(
        \i_fifo_rx/mem[35][5] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n484 ) );
  IMUX40 \i_fifo_rx/U520  ( .A(\i_fifo_rx/mem[36][5] ), .B(
        \i_fifo_rx/mem[37][5] ), .C(\i_fifo_rx/mem[38][5] ), .D(
        \i_fifo_rx/mem[39][5] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n486 ) );
  IMUX40 \i_fifo_rx/U420  ( .A(\i_fifo_rx/n484 ), .B(\i_fifo_rx/n485 ), .C(
        \i_fifo_rx/n486 ), .D(\i_fifo_rx/n487 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n483 ) );
  IMUX40 \i_fifo_rx/U515  ( .A(\i_fifo_rx/mem[56][5] ), .B(
        \i_fifo_rx/mem[57][5] ), .C(\i_fifo_rx/mem[58][5] ), .D(
        \i_fifo_rx/mem[59][5] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n480 ) );
  IMUX40 \i_fifo_rx/U517  ( .A(\i_fifo_rx/mem[48][5] ), .B(
        \i_fifo_rx/mem[49][5] ), .C(\i_fifo_rx/mem[50][5] ), .D(
        \i_fifo_rx/mem[51][5] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n479 ) );
  IMUX40 \i_fifo_rx/U516  ( .A(\i_fifo_rx/mem[52][5] ), .B(
        \i_fifo_rx/mem[53][5] ), .C(\i_fifo_rx/mem[54][5] ), .D(
        \i_fifo_rx/mem[55][5] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n481 ) );
  IMUX40 \i_fifo_rx/U419  ( .A(\i_fifo_rx/n479 ), .B(\i_fifo_rx/n480 ), .C(
        \i_fifo_rx/n481 ), .D(\i_fifo_rx/n482 ), .S0(\i_fifo_rx/N42 ), .S1(
        \i_fifo_rx/N41 ), .Q(\i_fifo_rx/n478 ) );
  IMUX40 \i_fifo_rx/U524  ( .A(\i_fifo_rx/mem[20][5] ), .B(
        \i_fifo_rx/mem[21][5] ), .C(\i_fifo_rx/mem[22][5] ), .D(
        \i_fifo_rx/mem[23][5] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n491 ) );
  IMUX40 \i_fifo_rx/U525  ( .A(\i_fifo_rx/mem[16][5] ), .B(
        \i_fifo_rx/mem[17][5] ), .C(\i_fifo_rx/mem[18][5] ), .D(
        \i_fifo_rx/mem[19][5] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n489 ) );
  IMUX40 \i_fifo_rx/U523  ( .A(\i_fifo_rx/mem[24][5] ), .B(
        \i_fifo_rx/mem[25][5] ), .C(\i_fifo_rx/mem[26][5] ), .D(
        \i_fifo_rx/mem[27][5] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n490 ) );
  IMUX40 \i_fifo_rx/U522  ( .A(\i_fifo_rx/mem[28][5] ), .B(
        \i_fifo_rx/mem[29][5] ), .C(\i_fifo_rx/mem[30][5] ), .D(
        \i_fifo_rx/mem[31][5] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n492 ) );
  IMUX40 \i_fifo_rx/U543  ( .A(\i_fifo_rx/mem[8][6] ), .B(
        \i_fifo_rx/mem[9][6] ), .C(\i_fifo_rx/mem[10][6] ), .D(
        \i_fifo_rx/mem[11][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n515 ) );
  IMUX40 \i_fifo_rx/U545  ( .A(\i_fifo_rx/mem[0][6] ), .B(
        \i_fifo_rx/mem[1][6] ), .C(\i_fifo_rx/mem[2][6] ), .D(
        \i_fifo_rx/mem[3][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n514 ) );
  IMUX40 \i_fifo_rx/U544  ( .A(\i_fifo_rx/mem[4][6] ), .B(
        \i_fifo_rx/mem[5][6] ), .C(\i_fifo_rx/mem[6][6] ), .D(
        \i_fifo_rx/mem[7][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n516 ) );
  IMUX40 \i_fifo_rx/U427  ( .A(\i_fifo_rx/n514 ), .B(\i_fifo_rx/n515 ), .C(
        \i_fifo_rx/n516 ), .D(\i_fifo_rx/n517 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n513 ) );
  IMUX40 \i_fifo_rx/U535  ( .A(\i_fifo_rx/mem[40][6] ), .B(
        \i_fifo_rx/mem[41][6] ), .C(\i_fifo_rx/mem[42][6] ), .D(
        \i_fifo_rx/mem[43][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n505 ) );
  IMUX40 \i_fifo_rx/U537  ( .A(\i_fifo_rx/mem[32][6] ), .B(
        \i_fifo_rx/mem[33][6] ), .C(\i_fifo_rx/mem[34][6] ), .D(
        \i_fifo_rx/mem[35][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n504 ) );
  IMUX40 \i_fifo_rx/U536  ( .A(\i_fifo_rx/mem[36][6] ), .B(
        \i_fifo_rx/mem[37][6] ), .C(\i_fifo_rx/mem[38][6] ), .D(
        \i_fifo_rx/mem[39][6] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n506 ) );
  IMUX40 \i_fifo_rx/U425  ( .A(\i_fifo_rx/n504 ), .B(\i_fifo_rx/n505 ), .C(
        \i_fifo_rx/n506 ), .D(\i_fifo_rx/n507 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n503 ) );
  IMUX40 \i_fifo_rx/U531  ( .A(\i_fifo_rx/mem[56][6] ), .B(
        \i_fifo_rx/mem[57][6] ), .C(\i_fifo_rx/mem[58][6] ), .D(
        \i_fifo_rx/mem[59][6] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n500 ) );
  IMUX40 \i_fifo_rx/U533  ( .A(\i_fifo_rx/mem[48][6] ), .B(
        \i_fifo_rx/mem[49][6] ), .C(\i_fifo_rx/mem[50][6] ), .D(
        \i_fifo_rx/mem[51][6] ), .S0(\i_fifo_rx/N39 ), .S1(n311), .Q(
        \i_fifo_rx/n499 ) );
  IMUX40 \i_fifo_rx/U532  ( .A(\i_fifo_rx/mem[52][6] ), .B(
        \i_fifo_rx/mem[53][6] ), .C(\i_fifo_rx/mem[54][6] ), .D(
        \i_fifo_rx/mem[55][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n501 ) );
  IMUX40 \i_fifo_rx/U424  ( .A(\i_fifo_rx/n499 ), .B(\i_fifo_rx/n500 ), .C(
        \i_fifo_rx/n501 ), .D(\i_fifo_rx/n502 ), .S0(\i_fifo_rx/N42 ), .S1(
        \i_fifo_rx/N41 ), .Q(\i_fifo_rx/n498 ) );
  IMUX40 \i_fifo_rx/U540  ( .A(\i_fifo_rx/mem[20][6] ), .B(
        \i_fifo_rx/mem[21][6] ), .C(\i_fifo_rx/mem[22][6] ), .D(
        \i_fifo_rx/mem[23][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n511 ) );
  IMUX40 \i_fifo_rx/U541  ( .A(\i_fifo_rx/mem[16][6] ), .B(
        \i_fifo_rx/mem[17][6] ), .C(\i_fifo_rx/mem[18][6] ), .D(
        \i_fifo_rx/mem[19][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n509 ) );
  IMUX40 \i_fifo_rx/U539  ( .A(\i_fifo_rx/mem[24][6] ), .B(
        \i_fifo_rx/mem[25][6] ), .C(\i_fifo_rx/mem[26][6] ), .D(
        \i_fifo_rx/mem[27][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n510 ) );
  IMUX40 \i_fifo_rx/U538  ( .A(\i_fifo_rx/mem[28][6] ), .B(
        \i_fifo_rx/mem[29][6] ), .C(\i_fifo_rx/mem[30][6] ), .D(
        \i_fifo_rx/mem[31][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n512 ) );
  IMUX40 \i_fifo_rx/U561  ( .A(\i_fifo_rx/mem[0][7] ), .B(
        \i_fifo_rx/mem[1][7] ), .C(\i_fifo_rx/mem[2][7] ), .D(
        \i_fifo_rx/mem[3][7] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n534 ) );
  IMUX40 \i_fifo_rx/U559  ( .A(\i_fifo_rx/mem[8][7] ), .B(
        \i_fifo_rx/mem[9][7] ), .C(\i_fifo_rx/mem[10][7] ), .D(
        \i_fifo_rx/mem[11][7] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n535 ) );
  IMUX40 \i_fifo_rx/U560  ( .A(\i_fifo_rx/mem[4][7] ), .B(
        \i_fifo_rx/mem[5][7] ), .C(\i_fifo_rx/mem[6][7] ), .D(
        \i_fifo_rx/mem[7][7] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n536 ) );
  IMUX40 \i_fifo_rx/U432  ( .A(\i_fifo_rx/n534 ), .B(\i_fifo_rx/n535 ), .C(
        \i_fifo_rx/n536 ), .D(\i_fifo_rx/n537 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n533 ) );
  IMUX40 \i_fifo_rx/U551  ( .A(\i_fifo_rx/mem[40][7] ), .B(
        \i_fifo_rx/mem[41][7] ), .C(\i_fifo_rx/mem[42][7] ), .D(
        \i_fifo_rx/mem[43][7] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n525 ) );
  IMUX40 \i_fifo_rx/U553  ( .A(\i_fifo_rx/mem[32][7] ), .B(
        \i_fifo_rx/mem[33][7] ), .C(\i_fifo_rx/mem[34][7] ), .D(
        \i_fifo_rx/mem[35][7] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n524 ) );
  IMUX40 \i_fifo_rx/U552  ( .A(\i_fifo_rx/mem[36][7] ), .B(
        \i_fifo_rx/mem[37][7] ), .C(\i_fifo_rx/mem[38][7] ), .D(
        \i_fifo_rx/mem[39][7] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n526 ) );
  IMUX40 \i_fifo_rx/U430  ( .A(\i_fifo_rx/n524 ), .B(\i_fifo_rx/n525 ), .C(
        \i_fifo_rx/n526 ), .D(\i_fifo_rx/n527 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n523 ) );
  IMUX40 \i_fifo_rx/U547  ( .A(\i_fifo_rx/mem[56][7] ), .B(
        \i_fifo_rx/mem[57][7] ), .C(\i_fifo_rx/mem[58][7] ), .D(
        \i_fifo_rx/mem[59][7] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n520 ) );
  IMUX40 \i_fifo_rx/U548  ( .A(\i_fifo_rx/mem[52][7] ), .B(
        \i_fifo_rx/mem[53][7] ), .C(\i_fifo_rx/mem[54][7] ), .D(
        \i_fifo_rx/mem[55][7] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n521 ) );
  IMUX40 \i_fifo_rx/U549  ( .A(\i_fifo_rx/mem[48][7] ), .B(
        \i_fifo_rx/mem[49][7] ), .C(\i_fifo_rx/mem[50][7] ), .D(
        \i_fifo_rx/mem[51][7] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n519 ) );
  IMUX40 \i_fifo_rx/U429  ( .A(\i_fifo_rx/n519 ), .B(\i_fifo_rx/n520 ), .C(
        \i_fifo_rx/n521 ), .D(\i_fifo_rx/n522 ), .S0(\i_fifo_rx/N42 ), .S1(
        \i_fifo_rx/N41 ), .Q(\i_fifo_rx/n518 ) );
  IMUX40 \i_fifo_rx/U556  ( .A(\i_fifo_rx/mem[20][7] ), .B(
        \i_fifo_rx/mem[21][7] ), .C(\i_fifo_rx/mem[22][7] ), .D(
        \i_fifo_rx/mem[23][7] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n531 ) );
  IMUX40 \i_fifo_rx/U557  ( .A(\i_fifo_rx/mem[16][7] ), .B(
        \i_fifo_rx/mem[17][7] ), .C(\i_fifo_rx/mem[18][7] ), .D(
        \i_fifo_rx/mem[19][7] ), .S0(n306), .S1(\i_fifo_rx/N40 ), .Q(
        \i_fifo_rx/n529 ) );
  IMUX40 \i_fifo_rx/U555  ( .A(\i_fifo_rx/mem[24][7] ), .B(
        \i_fifo_rx/mem[25][7] ), .C(\i_fifo_rx/mem[26][7] ), .D(
        \i_fifo_rx/mem[27][7] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n530 ) );
  IMUX40 \i_fifo_rx/U554  ( .A(\i_fifo_rx/mem[28][7] ), .B(
        \i_fifo_rx/mem[29][7] ), .C(\i_fifo_rx/mem[30][7] ), .D(
        \i_fifo_rx/mem[31][7] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n532 ) );
  IMUX40 \i_fifo_rx/U279  ( .A(\i_fifo_rx/mem[8][0] ), .B(
        \i_fifo_rx/mem[9][0] ), .C(\i_fifo_rx/mem[10][0] ), .D(
        \i_fifo_rx/mem[11][0] ), .S0(n302), .S1(n86), .Q(\i_fifo_rx/n235 ) );
  IMUX40 \i_fifo_rx/U281  ( .A(\i_fifo_rx/mem[0][0] ), .B(
        \i_fifo_rx/mem[1][0] ), .C(\i_fifo_rx/mem[2][0] ), .D(
        \i_fifo_rx/mem[3][0] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n234 ) );
  IMUX40 \i_fifo_rx/U280  ( .A(\i_fifo_rx/mem[4][0] ), .B(
        \i_fifo_rx/mem[5][0] ), .C(\i_fifo_rx/mem[6][0] ), .D(
        \i_fifo_rx/mem[7][0] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n236 ) );
  IMUX40 \i_fifo_rx/U229  ( .A(\i_fifo_rx/n234 ), .B(\i_fifo_rx/n235 ), .C(
        \i_fifo_rx/n236 ), .D(\i_fifo_rx/n237 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n233 ) );
  IMUX40 \i_fifo_rx/U271  ( .A(\i_fifo_rx/mem[40][0] ), .B(
        \i_fifo_rx/mem[41][0] ), .C(\i_fifo_rx/mem[42][0] ), .D(
        \i_fifo_rx/mem[43][0] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n225 ) );
  IMUX40 \i_fifo_rx/U273  ( .A(\i_fifo_rx/mem[32][0] ), .B(
        \i_fifo_rx/mem[33][0] ), .C(\i_fifo_rx/mem[34][0] ), .D(
        \i_fifo_rx/mem[35][0] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n224 ) );
  IMUX40 \i_fifo_rx/U272  ( .A(\i_fifo_rx/mem[36][0] ), .B(
        \i_fifo_rx/mem[37][0] ), .C(\i_fifo_rx/mem[38][0] ), .D(
        \i_fifo_rx/mem[39][0] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n226 ) );
  IMUX40 \i_fifo_rx/U227  ( .A(\i_fifo_rx/n224 ), .B(\i_fifo_rx/n225 ), .C(
        \i_fifo_rx/n226 ), .D(\i_fifo_rx/n227 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n223 ) );
  IMUX40 \i_fifo_rx/U267  ( .A(\i_fifo_rx/mem[56][0] ), .B(
        \i_fifo_rx/mem[57][0] ), .C(\i_fifo_rx/mem[58][0] ), .D(
        \i_fifo_rx/mem[59][0] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n220 ) );
  IMUX40 \i_fifo_rx/U269  ( .A(\i_fifo_rx/mem[48][0] ), .B(
        \i_fifo_rx/mem[49][0] ), .C(\i_fifo_rx/mem[50][0] ), .D(
        \i_fifo_rx/mem[51][0] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n219 ) );
  IMUX40 \i_fifo_rx/U268  ( .A(\i_fifo_rx/mem[52][0] ), .B(
        \i_fifo_rx/mem[53][0] ), .C(\i_fifo_rx/mem[54][0] ), .D(
        \i_fifo_rx/mem[55][0] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n221 ) );
  IMUX40 \i_fifo_rx/U226  ( .A(\i_fifo_rx/n219 ), .B(\i_fifo_rx/n220 ), .C(
        \i_fifo_rx/n221 ), .D(\i_fifo_rx/n222 ), .S0(\i_fifo_rx/N36 ), .S1(
        \i_fifo_rx/N35 ), .Q(\i_fifo_rx/n218 ) );
  IMUX40 \i_fifo_rx/U276  ( .A(\i_fifo_rx/mem[20][0] ), .B(
        \i_fifo_rx/mem[21][0] ), .C(\i_fifo_rx/mem[22][0] ), .D(
        \i_fifo_rx/mem[23][0] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n231 ) );
  IMUX40 \i_fifo_rx/U277  ( .A(\i_fifo_rx/mem[16][0] ), .B(
        \i_fifo_rx/mem[17][0] ), .C(\i_fifo_rx/mem[18][0] ), .D(
        \i_fifo_rx/mem[19][0] ), .S0(n302), .S1(n86), .Q(\i_fifo_rx/n229 ) );
  IMUX40 \i_fifo_rx/U275  ( .A(\i_fifo_rx/mem[24][0] ), .B(
        \i_fifo_rx/mem[25][0] ), .C(\i_fifo_rx/mem[26][0] ), .D(
        \i_fifo_rx/mem[27][0] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n230 ) );
  IMUX40 \i_fifo_rx/U274  ( .A(\i_fifo_rx/mem[28][0] ), .B(
        \i_fifo_rx/mem[29][0] ), .C(\i_fifo_rx/mem[30][0] ), .D(
        \i_fifo_rx/mem[31][0] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n232 ) );
  IMUX40 \i_fifo_rx/U295  ( .A(\i_fifo_rx/mem[8][1] ), .B(
        \i_fifo_rx/mem[9][1] ), .C(\i_fifo_rx/mem[10][1] ), .D(
        \i_fifo_rx/mem[11][1] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n255 ) );
  IMUX40 \i_fifo_rx/U297  ( .A(\i_fifo_rx/mem[0][1] ), .B(
        \i_fifo_rx/mem[1][1] ), .C(\i_fifo_rx/mem[2][1] ), .D(
        \i_fifo_rx/mem[3][1] ), .S0(n300), .S1(n86), .Q(\i_fifo_rx/n254 ) );
  IMUX40 \i_fifo_rx/U296  ( .A(\i_fifo_rx/mem[4][1] ), .B(
        \i_fifo_rx/mem[5][1] ), .C(\i_fifo_rx/mem[6][1] ), .D(
        \i_fifo_rx/mem[7][1] ), .S0(n302), .S1(n86), .Q(\i_fifo_rx/n256 ) );
  IMUX40 \i_fifo_rx/U234  ( .A(\i_fifo_rx/n254 ), .B(\i_fifo_rx/n255 ), .C(
        \i_fifo_rx/n256 ), .D(\i_fifo_rx/n257 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n253 ) );
  IMUX40 \i_fifo_rx/U287  ( .A(\i_fifo_rx/mem[40][1] ), .B(
        \i_fifo_rx/mem[41][1] ), .C(\i_fifo_rx/mem[42][1] ), .D(
        \i_fifo_rx/mem[43][1] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n245 ) );
  IMUX40 \i_fifo_rx/U289  ( .A(\i_fifo_rx/mem[32][1] ), .B(
        \i_fifo_rx/mem[33][1] ), .C(\i_fifo_rx/mem[34][1] ), .D(
        \i_fifo_rx/mem[35][1] ), .S0(n302), .S1(n86), .Q(\i_fifo_rx/n244 ) );
  IMUX40 \i_fifo_rx/U288  ( .A(\i_fifo_rx/mem[36][1] ), .B(
        \i_fifo_rx/mem[37][1] ), .C(\i_fifo_rx/mem[38][1] ), .D(
        \i_fifo_rx/mem[39][1] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n246 ) );
  IMUX40 \i_fifo_rx/U232  ( .A(\i_fifo_rx/n244 ), .B(\i_fifo_rx/n245 ), .C(
        \i_fifo_rx/n246 ), .D(\i_fifo_rx/n247 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n243 ) );
  IMUX40 \i_fifo_rx/U283  ( .A(\i_fifo_rx/mem[56][1] ), .B(
        \i_fifo_rx/mem[57][1] ), .C(\i_fifo_rx/mem[58][1] ), .D(
        \i_fifo_rx/mem[59][1] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n240 ) );
  IMUX40 \i_fifo_rx/U285  ( .A(\i_fifo_rx/mem[48][1] ), .B(
        \i_fifo_rx/mem[49][1] ), .C(\i_fifo_rx/mem[50][1] ), .D(
        \i_fifo_rx/mem[51][1] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n239 ) );
  IMUX40 \i_fifo_rx/U284  ( .A(\i_fifo_rx/mem[52][1] ), .B(
        \i_fifo_rx/mem[53][1] ), .C(\i_fifo_rx/mem[54][1] ), .D(
        \i_fifo_rx/mem[55][1] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n241 ) );
  IMUX40 \i_fifo_rx/U231  ( .A(\i_fifo_rx/n239 ), .B(\i_fifo_rx/n240 ), .C(
        \i_fifo_rx/n241 ), .D(\i_fifo_rx/n242 ), .S0(\i_fifo_rx/N36 ), .S1(
        n1945), .Q(\i_fifo_rx/n238 ) );
  IMUX40 \i_fifo_rx/U292  ( .A(\i_fifo_rx/mem[20][1] ), .B(
        \i_fifo_rx/mem[21][1] ), .C(\i_fifo_rx/mem[22][1] ), .D(
        \i_fifo_rx/mem[23][1] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n251 ) );
  IMUX40 \i_fifo_rx/U293  ( .A(\i_fifo_rx/mem[16][1] ), .B(
        \i_fifo_rx/mem[17][1] ), .C(\i_fifo_rx/mem[18][1] ), .D(
        \i_fifo_rx/mem[19][1] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n249 ) );
  IMUX40 \i_fifo_rx/U291  ( .A(\i_fifo_rx/mem[24][1] ), .B(
        \i_fifo_rx/mem[25][1] ), .C(\i_fifo_rx/mem[26][1] ), .D(
        \i_fifo_rx/mem[27][1] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n250 ) );
  IMUX40 \i_fifo_rx/U290  ( .A(\i_fifo_rx/mem[28][1] ), .B(
        \i_fifo_rx/mem[29][1] ), .C(\i_fifo_rx/mem[30][1] ), .D(
        \i_fifo_rx/mem[31][1] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n252 ) );
  IMUX40 \i_fifo_rx/U311  ( .A(\i_fifo_rx/mem[8][2] ), .B(
        \i_fifo_rx/mem[9][2] ), .C(\i_fifo_rx/mem[10][2] ), .D(
        \i_fifo_rx/mem[11][2] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n275 ) );
  IMUX40 \i_fifo_rx/U313  ( .A(\i_fifo_rx/mem[0][2] ), .B(
        \i_fifo_rx/mem[1][2] ), .C(\i_fifo_rx/mem[2][2] ), .D(
        \i_fifo_rx/mem[3][2] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n274 ) );
  IMUX40 \i_fifo_rx/U312  ( .A(\i_fifo_rx/mem[4][2] ), .B(
        \i_fifo_rx/mem[5][2] ), .C(\i_fifo_rx/mem[6][2] ), .D(
        \i_fifo_rx/mem[7][2] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n276 ) );
  IMUX40 \i_fifo_rx/U239  ( .A(\i_fifo_rx/n274 ), .B(\i_fifo_rx/n275 ), .C(
        \i_fifo_rx/n276 ), .D(\i_fifo_rx/n277 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n273 ) );
  IMUX40 \i_fifo_rx/U303  ( .A(\i_fifo_rx/mem[40][2] ), .B(
        \i_fifo_rx/mem[41][2] ), .C(\i_fifo_rx/mem[42][2] ), .D(
        \i_fifo_rx/mem[43][2] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n265 ) );
  IMUX40 \i_fifo_rx/U305  ( .A(\i_fifo_rx/mem[32][2] ), .B(
        \i_fifo_rx/mem[33][2] ), .C(\i_fifo_rx/mem[34][2] ), .D(
        \i_fifo_rx/mem[35][2] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n264 ) );
  IMUX40 \i_fifo_rx/U304  ( .A(\i_fifo_rx/mem[36][2] ), .B(
        \i_fifo_rx/mem[37][2] ), .C(\i_fifo_rx/mem[38][2] ), .D(
        \i_fifo_rx/mem[39][2] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n266 ) );
  IMUX40 \i_fifo_rx/U237  ( .A(\i_fifo_rx/n264 ), .B(\i_fifo_rx/n265 ), .C(
        \i_fifo_rx/n266 ), .D(\i_fifo_rx/n267 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n263 ) );
  IMUX40 \i_fifo_rx/U299  ( .A(\i_fifo_rx/mem[56][2] ), .B(
        \i_fifo_rx/mem[57][2] ), .C(\i_fifo_rx/mem[58][2] ), .D(
        \i_fifo_rx/mem[59][2] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n260 ) );
  IMUX40 \i_fifo_rx/U301  ( .A(\i_fifo_rx/mem[48][2] ), .B(
        \i_fifo_rx/mem[49][2] ), .C(\i_fifo_rx/mem[50][2] ), .D(
        \i_fifo_rx/mem[51][2] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n259 ) );
  IMUX40 \i_fifo_rx/U300  ( .A(\i_fifo_rx/mem[52][2] ), .B(
        \i_fifo_rx/mem[53][2] ), .C(\i_fifo_rx/mem[54][2] ), .D(
        \i_fifo_rx/mem[55][2] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n261 ) );
  IMUX40 \i_fifo_rx/U236  ( .A(\i_fifo_rx/n259 ), .B(\i_fifo_rx/n260 ), .C(
        \i_fifo_rx/n261 ), .D(\i_fifo_rx/n262 ), .S0(\i_fifo_rx/N36 ), .S1(
        \i_fifo_rx/N35 ), .Q(\i_fifo_rx/n258 ) );
  IMUX40 \i_fifo_rx/U308  ( .A(\i_fifo_rx/mem[20][2] ), .B(
        \i_fifo_rx/mem[21][2] ), .C(\i_fifo_rx/mem[22][2] ), .D(
        \i_fifo_rx/mem[23][2] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n271 ) );
  IMUX40 \i_fifo_rx/U309  ( .A(\i_fifo_rx/mem[16][2] ), .B(
        \i_fifo_rx/mem[17][2] ), .C(\i_fifo_rx/mem[18][2] ), .D(
        \i_fifo_rx/mem[19][2] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n269 ) );
  IMUX40 \i_fifo_rx/U307  ( .A(\i_fifo_rx/mem[24][2] ), .B(
        \i_fifo_rx/mem[25][2] ), .C(\i_fifo_rx/mem[26][2] ), .D(
        \i_fifo_rx/mem[27][2] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n270 ) );
  IMUX40 \i_fifo_rx/U306  ( .A(\i_fifo_rx/mem[28][2] ), .B(
        \i_fifo_rx/mem[29][2] ), .C(\i_fifo_rx/mem[30][2] ), .D(
        \i_fifo_rx/mem[31][2] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n272 ) );
  IMUX40 \i_fifo_rx/U327  ( .A(\i_fifo_rx/mem[8][3] ), .B(
        \i_fifo_rx/mem[9][3] ), .C(\i_fifo_rx/mem[10][3] ), .D(
        \i_fifo_rx/mem[11][3] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n295 ) );
  IMUX40 \i_fifo_rx/U329  ( .A(\i_fifo_rx/mem[0][3] ), .B(
        \i_fifo_rx/mem[1][3] ), .C(\i_fifo_rx/mem[2][3] ), .D(
        \i_fifo_rx/mem[3][3] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n294 ) );
  IMUX40 \i_fifo_rx/U328  ( .A(\i_fifo_rx/mem[4][3] ), .B(
        \i_fifo_rx/mem[5][3] ), .C(\i_fifo_rx/mem[6][3] ), .D(
        \i_fifo_rx/mem[7][3] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n296 ) );
  IMUX40 \i_fifo_rx/U244  ( .A(\i_fifo_rx/n294 ), .B(\i_fifo_rx/n295 ), .C(
        \i_fifo_rx/n296 ), .D(\i_fifo_rx/n297 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n293 ) );
  IMUX40 \i_fifo_rx/U319  ( .A(\i_fifo_rx/mem[40][3] ), .B(
        \i_fifo_rx/mem[41][3] ), .C(\i_fifo_rx/mem[42][3] ), .D(
        \i_fifo_rx/mem[43][3] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n285 ) );
  IMUX40 \i_fifo_rx/U321  ( .A(\i_fifo_rx/mem[32][3] ), .B(
        \i_fifo_rx/mem[33][3] ), .C(\i_fifo_rx/mem[34][3] ), .D(
        \i_fifo_rx/mem[35][3] ), .S0(n300), .S1(n86), .Q(\i_fifo_rx/n284 ) );
  IMUX40 \i_fifo_rx/U320  ( .A(\i_fifo_rx/mem[36][3] ), .B(
        \i_fifo_rx/mem[37][3] ), .C(\i_fifo_rx/mem[38][3] ), .D(
        \i_fifo_rx/mem[39][3] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n286 ) );
  IMUX40 \i_fifo_rx/U242  ( .A(\i_fifo_rx/n284 ), .B(\i_fifo_rx/n285 ), .C(
        \i_fifo_rx/n286 ), .D(\i_fifo_rx/n287 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n283 ) );
  IMUX40 \i_fifo_rx/U315  ( .A(\i_fifo_rx/mem[56][3] ), .B(
        \i_fifo_rx/mem[57][3] ), .C(\i_fifo_rx/mem[58][3] ), .D(
        \i_fifo_rx/mem[59][3] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n280 ) );
  IMUX40 \i_fifo_rx/U317  ( .A(\i_fifo_rx/mem[48][3] ), .B(
        \i_fifo_rx/mem[49][3] ), .C(\i_fifo_rx/mem[50][3] ), .D(
        \i_fifo_rx/mem[51][3] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n279 ) );
  IMUX40 \i_fifo_rx/U316  ( .A(\i_fifo_rx/mem[52][3] ), .B(
        \i_fifo_rx/mem[53][3] ), .C(\i_fifo_rx/mem[54][3] ), .D(
        \i_fifo_rx/mem[55][3] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n281 ) );
  IMUX40 \i_fifo_rx/U241  ( .A(\i_fifo_rx/n279 ), .B(\i_fifo_rx/n280 ), .C(
        \i_fifo_rx/n281 ), .D(\i_fifo_rx/n282 ), .S0(\i_fifo_rx/N36 ), .S1(
        \i_fifo_rx/N35 ), .Q(\i_fifo_rx/n278 ) );
  IMUX40 \i_fifo_rx/U324  ( .A(\i_fifo_rx/mem[20][3] ), .B(
        \i_fifo_rx/mem[21][3] ), .C(\i_fifo_rx/mem[22][3] ), .D(
        \i_fifo_rx/mem[23][3] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n291 ) );
  IMUX40 \i_fifo_rx/U325  ( .A(\i_fifo_rx/mem[16][3] ), .B(
        \i_fifo_rx/mem[17][3] ), .C(\i_fifo_rx/mem[18][3] ), .D(
        \i_fifo_rx/mem[19][3] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n289 ) );
  IMUX40 \i_fifo_rx/U323  ( .A(\i_fifo_rx/mem[24][3] ), .B(
        \i_fifo_rx/mem[25][3] ), .C(\i_fifo_rx/mem[26][3] ), .D(
        \i_fifo_rx/mem[27][3] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n290 ) );
  IMUX40 \i_fifo_rx/U322  ( .A(\i_fifo_rx/mem[28][3] ), .B(
        \i_fifo_rx/mem[29][3] ), .C(\i_fifo_rx/mem[30][3] ), .D(
        \i_fifo_rx/mem[31][3] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n292 ) );
  IMUX40 \i_fifo_rx/U343  ( .A(\i_fifo_rx/mem[8][4] ), .B(
        \i_fifo_rx/mem[9][4] ), .C(\i_fifo_rx/mem[10][4] ), .D(
        \i_fifo_rx/mem[11][4] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n315 ) );
  IMUX40 \i_fifo_rx/U345  ( .A(\i_fifo_rx/mem[0][4] ), .B(
        \i_fifo_rx/mem[1][4] ), .C(\i_fifo_rx/mem[2][4] ), .D(
        \i_fifo_rx/mem[3][4] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n314 ) );
  IMUX40 \i_fifo_rx/U344  ( .A(\i_fifo_rx/mem[4][4] ), .B(
        \i_fifo_rx/mem[5][4] ), .C(\i_fifo_rx/mem[6][4] ), .D(
        \i_fifo_rx/mem[7][4] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n316 ) );
  IMUX40 \i_fifo_rx/U249  ( .A(\i_fifo_rx/n314 ), .B(\i_fifo_rx/n315 ), .C(
        \i_fifo_rx/n316 ), .D(\i_fifo_rx/n317 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n313 ) );
  IMUX40 \i_fifo_rx/U335  ( .A(\i_fifo_rx/mem[40][4] ), .B(
        \i_fifo_rx/mem[41][4] ), .C(\i_fifo_rx/mem[42][4] ), .D(
        \i_fifo_rx/mem[43][4] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n305 ) );
  IMUX40 \i_fifo_rx/U337  ( .A(\i_fifo_rx/mem[32][4] ), .B(
        \i_fifo_rx/mem[33][4] ), .C(\i_fifo_rx/mem[34][4] ), .D(
        \i_fifo_rx/mem[35][4] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n304 ) );
  IMUX40 \i_fifo_rx/U336  ( .A(\i_fifo_rx/mem[36][4] ), .B(
        \i_fifo_rx/mem[37][4] ), .C(\i_fifo_rx/mem[38][4] ), .D(
        \i_fifo_rx/mem[39][4] ), .S0(n134), .S1(n305), .Q(\i_fifo_rx/n306 ) );
  IMUX40 \i_fifo_rx/U247  ( .A(\i_fifo_rx/n304 ), .B(\i_fifo_rx/n305 ), .C(
        \i_fifo_rx/n306 ), .D(\i_fifo_rx/n307 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n303 ) );
  IMUX40 \i_fifo_rx/U331  ( .A(\i_fifo_rx/mem[56][4] ), .B(
        \i_fifo_rx/mem[57][4] ), .C(\i_fifo_rx/mem[58][4] ), .D(
        \i_fifo_rx/mem[59][4] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n300 ) );
  IMUX40 \i_fifo_rx/U333  ( .A(\i_fifo_rx/mem[48][4] ), .B(
        \i_fifo_rx/mem[49][4] ), .C(\i_fifo_rx/mem[50][4] ), .D(
        \i_fifo_rx/mem[51][4] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n299 ) );
  IMUX40 \i_fifo_rx/U332  ( .A(\i_fifo_rx/mem[52][4] ), .B(
        \i_fifo_rx/mem[53][4] ), .C(\i_fifo_rx/mem[54][4] ), .D(
        \i_fifo_rx/mem[55][4] ), .S0(n134), .S1(n305), .Q(\i_fifo_rx/n301 ) );
  IMUX40 \i_fifo_rx/U246  ( .A(\i_fifo_rx/n299 ), .B(\i_fifo_rx/n300 ), .C(
        \i_fifo_rx/n301 ), .D(\i_fifo_rx/n302 ), .S0(\i_fifo_rx/N36 ), .S1(
        \i_fifo_rx/N35 ), .Q(\i_fifo_rx/n298 ) );
  IMUX40 \i_fifo_rx/U340  ( .A(\i_fifo_rx/mem[20][4] ), .B(
        \i_fifo_rx/mem[21][4] ), .C(\i_fifo_rx/mem[22][4] ), .D(
        \i_fifo_rx/mem[23][4] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n311 ) );
  IMUX40 \i_fifo_rx/U341  ( .A(\i_fifo_rx/mem[16][4] ), .B(
        \i_fifo_rx/mem[17][4] ), .C(\i_fifo_rx/mem[18][4] ), .D(
        \i_fifo_rx/mem[19][4] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n309 ) );
  IMUX40 \i_fifo_rx/U339  ( .A(\i_fifo_rx/mem[24][4] ), .B(
        \i_fifo_rx/mem[25][4] ), .C(\i_fifo_rx/mem[26][4] ), .D(
        \i_fifo_rx/mem[27][4] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n310 ) );
  IMUX40 \i_fifo_rx/U338  ( .A(\i_fifo_rx/mem[28][4] ), .B(
        \i_fifo_rx/mem[29][4] ), .C(\i_fifo_rx/mem[30][4] ), .D(
        \i_fifo_rx/mem[31][4] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n312 ) );
  IMUX40 \i_fifo_rx/U359  ( .A(\i_fifo_rx/mem[8][5] ), .B(
        \i_fifo_rx/mem[9][5] ), .C(\i_fifo_rx/mem[10][5] ), .D(
        \i_fifo_rx/mem[11][5] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n335 ) );
  IMUX40 \i_fifo_rx/U361  ( .A(\i_fifo_rx/mem[0][5] ), .B(
        \i_fifo_rx/mem[1][5] ), .C(\i_fifo_rx/mem[2][5] ), .D(
        \i_fifo_rx/mem[3][5] ), .S0(n300), .S1(n86), .Q(\i_fifo_rx/n334 ) );
  IMUX40 \i_fifo_rx/U360  ( .A(\i_fifo_rx/mem[4][5] ), .B(
        \i_fifo_rx/mem[5][5] ), .C(\i_fifo_rx/mem[6][5] ), .D(
        \i_fifo_rx/mem[7][5] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n336 ) );
  IMUX40 \i_fifo_rx/U254  ( .A(\i_fifo_rx/n334 ), .B(\i_fifo_rx/n335 ), .C(
        \i_fifo_rx/n336 ), .D(\i_fifo_rx/n337 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n333 ) );
  IMUX40 \i_fifo_rx/U351  ( .A(\i_fifo_rx/mem[40][5] ), .B(
        \i_fifo_rx/mem[41][5] ), .C(\i_fifo_rx/mem[42][5] ), .D(
        \i_fifo_rx/mem[43][5] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n325 ) );
  IMUX40 \i_fifo_rx/U353  ( .A(\i_fifo_rx/mem[32][5] ), .B(
        \i_fifo_rx/mem[33][5] ), .C(\i_fifo_rx/mem[34][5] ), .D(
        \i_fifo_rx/mem[35][5] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n324 ) );
  IMUX40 \i_fifo_rx/U352  ( .A(\i_fifo_rx/mem[36][5] ), .B(
        \i_fifo_rx/mem[37][5] ), .C(\i_fifo_rx/mem[38][5] ), .D(
        \i_fifo_rx/mem[39][5] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n326 ) );
  IMUX40 \i_fifo_rx/U252  ( .A(\i_fifo_rx/n324 ), .B(\i_fifo_rx/n325 ), .C(
        \i_fifo_rx/n326 ), .D(\i_fifo_rx/n327 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n323 ) );
  IMUX40 \i_fifo_rx/U347  ( .A(\i_fifo_rx/mem[56][5] ), .B(
        \i_fifo_rx/mem[57][5] ), .C(\i_fifo_rx/mem[58][5] ), .D(
        \i_fifo_rx/mem[59][5] ), .S0(n134), .S1(n305), .Q(\i_fifo_rx/n320 ) );
  IMUX40 \i_fifo_rx/U349  ( .A(\i_fifo_rx/mem[48][5] ), .B(
        \i_fifo_rx/mem[49][5] ), .C(\i_fifo_rx/mem[50][5] ), .D(
        \i_fifo_rx/mem[51][5] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n319 ) );
  IMUX40 \i_fifo_rx/U348  ( .A(\i_fifo_rx/mem[52][5] ), .B(
        \i_fifo_rx/mem[53][5] ), .C(\i_fifo_rx/mem[54][5] ), .D(
        \i_fifo_rx/mem[55][5] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n321 ) );
  IMUX40 \i_fifo_rx/U251  ( .A(\i_fifo_rx/n319 ), .B(\i_fifo_rx/n320 ), .C(
        \i_fifo_rx/n321 ), .D(\i_fifo_rx/n322 ), .S0(\i_fifo_rx/N36 ), .S1(
        n1945), .Q(\i_fifo_rx/n318 ) );
  IMUX40 \i_fifo_rx/U356  ( .A(\i_fifo_rx/mem[20][5] ), .B(
        \i_fifo_rx/mem[21][5] ), .C(\i_fifo_rx/mem[22][5] ), .D(
        \i_fifo_rx/mem[23][5] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n331 ) );
  IMUX40 \i_fifo_rx/U357  ( .A(\i_fifo_rx/mem[16][5] ), .B(
        \i_fifo_rx/mem[17][5] ), .C(\i_fifo_rx/mem[18][5] ), .D(
        \i_fifo_rx/mem[19][5] ), .S0(n300), .S1(n86), .Q(\i_fifo_rx/n329 ) );
  IMUX40 \i_fifo_rx/U355  ( .A(\i_fifo_rx/mem[24][5] ), .B(
        \i_fifo_rx/mem[25][5] ), .C(\i_fifo_rx/mem[26][5] ), .D(
        \i_fifo_rx/mem[27][5] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n330 ) );
  IMUX40 \i_fifo_rx/U354  ( .A(\i_fifo_rx/mem[28][5] ), .B(
        \i_fifo_rx/mem[29][5] ), .C(\i_fifo_rx/mem[30][5] ), .D(
        \i_fifo_rx/mem[31][5] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n332 ) );
  IMUX40 \i_fifo_rx/U375  ( .A(\i_fifo_rx/mem[8][6] ), .B(
        \i_fifo_rx/mem[9][6] ), .C(\i_fifo_rx/mem[10][6] ), .D(
        \i_fifo_rx/mem[11][6] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n355 ) );
  IMUX40 \i_fifo_rx/U377  ( .A(\i_fifo_rx/mem[0][6] ), .B(
        \i_fifo_rx/mem[1][6] ), .C(\i_fifo_rx/mem[2][6] ), .D(
        \i_fifo_rx/mem[3][6] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n354 ) );
  IMUX40 \i_fifo_rx/U376  ( .A(\i_fifo_rx/mem[4][6] ), .B(
        \i_fifo_rx/mem[5][6] ), .C(\i_fifo_rx/mem[6][6] ), .D(
        \i_fifo_rx/mem[7][6] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n356 ) );
  IMUX40 \i_fifo_rx/U259  ( .A(\i_fifo_rx/n354 ), .B(\i_fifo_rx/n355 ), .C(
        \i_fifo_rx/n356 ), .D(\i_fifo_rx/n357 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n353 ) );
  IMUX40 \i_fifo_rx/U367  ( .A(\i_fifo_rx/mem[40][6] ), .B(
        \i_fifo_rx/mem[41][6] ), .C(\i_fifo_rx/mem[42][6] ), .D(
        \i_fifo_rx/mem[43][6] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n345 ) );
  IMUX40 \i_fifo_rx/U368  ( .A(\i_fifo_rx/mem[36][6] ), .B(
        \i_fifo_rx/mem[37][6] ), .C(\i_fifo_rx/mem[38][6] ), .D(
        \i_fifo_rx/mem[39][6] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n346 ) );
  IMUX40 \i_fifo_rx/U369  ( .A(\i_fifo_rx/mem[32][6] ), .B(
        \i_fifo_rx/mem[33][6] ), .C(\i_fifo_rx/mem[34][6] ), .D(
        \i_fifo_rx/mem[35][6] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n344 ) );
  IMUX40 \i_fifo_rx/U257  ( .A(\i_fifo_rx/n344 ), .B(\i_fifo_rx/n345 ), .C(
        \i_fifo_rx/n346 ), .D(\i_fifo_rx/n347 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n343 ) );
  IMUX40 \i_fifo_rx/U363  ( .A(\i_fifo_rx/mem[56][6] ), .B(
        \i_fifo_rx/mem[57][6] ), .C(\i_fifo_rx/mem[58][6] ), .D(
        \i_fifo_rx/mem[59][6] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n340 ) );
  IMUX40 \i_fifo_rx/U365  ( .A(\i_fifo_rx/mem[48][6] ), .B(
        \i_fifo_rx/mem[49][6] ), .C(\i_fifo_rx/mem[50][6] ), .D(
        \i_fifo_rx/mem[51][6] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n339 ) );
  IMUX40 \i_fifo_rx/U364  ( .A(\i_fifo_rx/mem[52][6] ), .B(
        \i_fifo_rx/mem[53][6] ), .C(\i_fifo_rx/mem[54][6] ), .D(
        \i_fifo_rx/mem[55][6] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n341 ) );
  IMUX40 \i_fifo_rx/U256  ( .A(\i_fifo_rx/n339 ), .B(\i_fifo_rx/n340 ), .C(
        \i_fifo_rx/n341 ), .D(\i_fifo_rx/n342 ), .S0(\i_fifo_rx/N36 ), .S1(
        n1945), .Q(\i_fifo_rx/n338 ) );
  IMUX40 \i_fifo_rx/U372  ( .A(\i_fifo_rx/mem[20][6] ), .B(
        \i_fifo_rx/mem[21][6] ), .C(\i_fifo_rx/mem[22][6] ), .D(
        \i_fifo_rx/mem[23][6] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n351 ) );
  IMUX40 \i_fifo_rx/U373  ( .A(\i_fifo_rx/mem[16][6] ), .B(
        \i_fifo_rx/mem[17][6] ), .C(\i_fifo_rx/mem[18][6] ), .D(
        \i_fifo_rx/mem[19][6] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n349 ) );
  IMUX40 \i_fifo_rx/U371  ( .A(\i_fifo_rx/mem[24][6] ), .B(
        \i_fifo_rx/mem[25][6] ), .C(\i_fifo_rx/mem[26][6] ), .D(
        \i_fifo_rx/mem[27][6] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n350 ) );
  IMUX40 \i_fifo_rx/U370  ( .A(\i_fifo_rx/mem[28][6] ), .B(
        \i_fifo_rx/mem[29][6] ), .C(\i_fifo_rx/mem[30][6] ), .D(
        \i_fifo_rx/mem[31][6] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n352 ) );
  IMUX40 \i_fifo_rx/U390  ( .A(\i_fifo_rx/mem[12][7] ), .B(
        \i_fifo_rx/mem[13][7] ), .C(\i_fifo_rx/mem[14][7] ), .D(
        \i_fifo_rx/mem[15][7] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n377 ) );
  IMUX40 \i_fifo_rx/U391  ( .A(\i_fifo_rx/mem[8][7] ), .B(
        \i_fifo_rx/mem[9][7] ), .C(\i_fifo_rx/mem[10][7] ), .D(
        \i_fifo_rx/mem[11][7] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n375 ) );
  IMUX40 \i_fifo_rx/U392  ( .A(\i_fifo_rx/mem[4][7] ), .B(
        \i_fifo_rx/mem[5][7] ), .C(\i_fifo_rx/mem[6][7] ), .D(
        \i_fifo_rx/mem[7][7] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n376 ) );
  IMUX40 \i_fifo_rx/U264  ( .A(\i_fifo_rx/n374 ), .B(\i_fifo_rx/n375 ), .C(
        \i_fifo_rx/n376 ), .D(\i_fifo_rx/n377 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n373 ) );
  IMUX40 \i_fifo_rx/U383  ( .A(\i_fifo_rx/mem[40][7] ), .B(
        \i_fifo_rx/mem[41][7] ), .C(\i_fifo_rx/mem[42][7] ), .D(
        \i_fifo_rx/mem[43][7] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n365 ) );
  IMUX40 \i_fifo_rx/U385  ( .A(\i_fifo_rx/mem[32][7] ), .B(
        \i_fifo_rx/mem[33][7] ), .C(\i_fifo_rx/mem[34][7] ), .D(
        \i_fifo_rx/mem[35][7] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n364 ) );
  IMUX40 \i_fifo_rx/U384  ( .A(\i_fifo_rx/mem[36][7] ), .B(
        \i_fifo_rx/mem[37][7] ), .C(\i_fifo_rx/mem[38][7] ), .D(
        \i_fifo_rx/mem[39][7] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n366 ) );
  IMUX40 \i_fifo_rx/U262  ( .A(\i_fifo_rx/n364 ), .B(\i_fifo_rx/n365 ), .C(
        \i_fifo_rx/n366 ), .D(\i_fifo_rx/n367 ), .S0(n274), .S1(n1945), .Q(
        \i_fifo_rx/n363 ) );
  IMUX40 \i_fifo_rx/U379  ( .A(\i_fifo_rx/mem[56][7] ), .B(
        \i_fifo_rx/mem[57][7] ), .C(\i_fifo_rx/mem[58][7] ), .D(
        \i_fifo_rx/mem[59][7] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n360 ) );
  IMUX40 \i_fifo_rx/U381  ( .A(\i_fifo_rx/mem[48][7] ), .B(
        \i_fifo_rx/mem[49][7] ), .C(\i_fifo_rx/mem[50][7] ), .D(
        \i_fifo_rx/mem[51][7] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n359 ) );
  IMUX40 \i_fifo_rx/U380  ( .A(\i_fifo_rx/mem[52][7] ), .B(
        \i_fifo_rx/mem[53][7] ), .C(\i_fifo_rx/mem[54][7] ), .D(
        \i_fifo_rx/mem[55][7] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n361 ) );
  IMUX40 \i_fifo_rx/U261  ( .A(\i_fifo_rx/n359 ), .B(\i_fifo_rx/n360 ), .C(
        \i_fifo_rx/n361 ), .D(\i_fifo_rx/n362 ), .S0(\i_fifo_rx/N36 ), .S1(
        n1945), .Q(\i_fifo_rx/n358 ) );
  IMUX40 \i_fifo_rx/U388  ( .A(\i_fifo_rx/mem[20][7] ), .B(
        \i_fifo_rx/mem[21][7] ), .C(\i_fifo_rx/mem[22][7] ), .D(
        \i_fifo_rx/mem[23][7] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n371 ) );
  IMUX40 \i_fifo_rx/U389  ( .A(\i_fifo_rx/mem[16][7] ), .B(
        \i_fifo_rx/mem[17][7] ), .C(\i_fifo_rx/mem[18][7] ), .D(
        \i_fifo_rx/mem[19][7] ), .S0(n299), .S1(n86), .Q(\i_fifo_rx/n369 ) );
  IMUX40 \i_fifo_rx/U387  ( .A(\i_fifo_rx/mem[24][7] ), .B(
        \i_fifo_rx/mem[25][7] ), .C(\i_fifo_rx/mem[26][7] ), .D(
        \i_fifo_rx/mem[27][7] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n370 ) );
  IMUX40 \i_fifo_rx/U386  ( .A(\i_fifo_rx/mem[28][7] ), .B(
        \i_fifo_rx/mem[29][7] ), .C(\i_fifo_rx/mem[30][7] ), .D(
        \i_fifo_rx/mem[31][7] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n372 ) );
  IMUX21 \i_fifo_tx/U542  ( .A(\i_fifo_tx/n528 ), .B(\i_fifo_tx/n529 ), .S(
        \i_fifo_tx/N38 ), .Q(\i_fifo_tx/N144 ) );
  IMUX40 \i_fifo_tx/U254  ( .A(\i_fifo_tx/mem[28][0] ), .B(
        \i_fifo_tx/mem[29][0] ), .C(\i_fifo_tx/mem[30][0] ), .D(
        \i_fifo_tx/mem[31][0] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n222 ) );
  IMUX40 \i_fifo_tx/U258  ( .A(\i_fifo_tx/mem[12][0] ), .B(
        \i_fifo_tx/mem[13][0] ), .C(\i_fifo_tx/mem[14][0] ), .D(
        \i_fifo_tx/mem[15][0] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n227 ) );
  IMUX40 \i_fifo_tx/U250  ( .A(\i_fifo_tx/mem[44][0] ), .B(
        \i_fifo_tx/mem[45][0] ), .C(\i_fifo_tx/mem[46][0] ), .D(
        \i_fifo_tx/mem[47][0] ), .S0(n317), .S1(n319), .Q(\i_fifo_tx/n217 ) );
  IMUX40 \i_fifo_tx/U246  ( .A(\i_fifo_tx/mem[60][0] ), .B(
        \i_fifo_tx/mem[61][0] ), .C(\i_fifo_tx/mem[62][0] ), .D(
        \i_fifo_tx/mem[63][0] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n212 ) );
  IMUX40 \i_fifo_tx/U270  ( .A(\i_fifo_tx/mem[28][1] ), .B(
        \i_fifo_tx/mem[29][1] ), .C(\i_fifo_tx/mem[30][1] ), .D(
        \i_fifo_tx/mem[31][1] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n242 ) );
  IMUX40 \i_fifo_tx/U274  ( .A(\i_fifo_tx/mem[12][1] ), .B(
        \i_fifo_tx/mem[13][1] ), .C(\i_fifo_tx/mem[14][1] ), .D(
        \i_fifo_tx/mem[15][1] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n247 ) );
  IMUX40 \i_fifo_tx/U266  ( .A(\i_fifo_tx/mem[44][1] ), .B(
        \i_fifo_tx/mem[45][1] ), .C(\i_fifo_tx/mem[46][1] ), .D(
        \i_fifo_tx/mem[47][1] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n237 ) );
  IMUX40 \i_fifo_tx/U262  ( .A(\i_fifo_tx/mem[60][1] ), .B(
        \i_fifo_tx/mem[61][1] ), .C(\i_fifo_tx/mem[62][1] ), .D(
        \i_fifo_tx/mem[63][1] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n232 ) );
  IMUX40 \i_fifo_tx/U286  ( .A(\i_fifo_tx/mem[28][2] ), .B(
        \i_fifo_tx/mem[29][2] ), .C(\i_fifo_tx/mem[30][2] ), .D(
        \i_fifo_tx/mem[31][2] ), .S0(n132), .S1(n318), .Q(\i_fifo_tx/n262 ) );
  IMUX40 \i_fifo_tx/U290  ( .A(\i_fifo_tx/mem[12][2] ), .B(
        \i_fifo_tx/mem[13][2] ), .C(\i_fifo_tx/mem[14][2] ), .D(
        \i_fifo_tx/mem[15][2] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n267 ) );
  IMUX40 \i_fifo_tx/U282  ( .A(\i_fifo_tx/mem[44][2] ), .B(
        \i_fifo_tx/mem[45][2] ), .C(\i_fifo_tx/mem[46][2] ), .D(
        \i_fifo_tx/mem[47][2] ), .S0(n132), .S1(n319), .Q(\i_fifo_tx/n257 ) );
  IMUX40 \i_fifo_tx/U278  ( .A(\i_fifo_tx/mem[60][2] ), .B(
        \i_fifo_tx/mem[61][2] ), .C(\i_fifo_tx/mem[62][2] ), .D(
        \i_fifo_tx/mem[63][2] ), .S0(n132), .S1(n318), .Q(\i_fifo_tx/n252 ) );
  IMUX40 \i_fifo_tx/U302  ( .A(\i_fifo_tx/mem[28][3] ), .B(
        \i_fifo_tx/mem[29][3] ), .C(\i_fifo_tx/mem[30][3] ), .D(
        \i_fifo_tx/mem[31][3] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n282 ) );
  IMUX40 \i_fifo_tx/U306  ( .A(\i_fifo_tx/mem[12][3] ), .B(
        \i_fifo_tx/mem[13][3] ), .C(\i_fifo_tx/mem[14][3] ), .D(
        \i_fifo_tx/mem[15][3] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n287 ) );
  IMUX40 \i_fifo_tx/U298  ( .A(\i_fifo_tx/mem[44][3] ), .B(
        \i_fifo_tx/mem[45][3] ), .C(\i_fifo_tx/mem[46][3] ), .D(
        \i_fifo_tx/mem[47][3] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n277 ) );
  IMUX40 \i_fifo_tx/U294  ( .A(\i_fifo_tx/mem[60][3] ), .B(
        \i_fifo_tx/mem[61][3] ), .C(\i_fifo_tx/mem[62][3] ), .D(
        \i_fifo_tx/mem[63][3] ), .S0(n316), .S1(n319), .Q(\i_fifo_tx/n272 ) );
  IMUX40 \i_fifo_tx/U318  ( .A(\i_fifo_tx/mem[28][4] ), .B(
        \i_fifo_tx/mem[29][4] ), .C(\i_fifo_tx/mem[30][4] ), .D(
        \i_fifo_tx/mem[31][4] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n302 ) );
  IMUX40 \i_fifo_tx/U322  ( .A(\i_fifo_tx/mem[12][4] ), .B(
        \i_fifo_tx/mem[13][4] ), .C(\i_fifo_tx/mem[14][4] ), .D(
        \i_fifo_tx/mem[15][4] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n307 ) );
  IMUX40 \i_fifo_tx/U314  ( .A(\i_fifo_tx/mem[44][4] ), .B(
        \i_fifo_tx/mem[45][4] ), .C(\i_fifo_tx/mem[46][4] ), .D(
        \i_fifo_tx/mem[47][4] ), .S0(n132), .S1(n318), .Q(\i_fifo_tx/n297 ) );
  IMUX40 \i_fifo_tx/U310  ( .A(\i_fifo_tx/mem[60][4] ), .B(
        \i_fifo_tx/mem[61][4] ), .C(\i_fifo_tx/mem[62][4] ), .D(
        \i_fifo_tx/mem[63][4] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n292 ) );
  IMUX40 \i_fifo_tx/U334  ( .A(\i_fifo_tx/mem[28][5] ), .B(
        \i_fifo_tx/mem[29][5] ), .C(\i_fifo_tx/mem[30][5] ), .D(
        \i_fifo_tx/mem[31][5] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n322 ) );
  IMUX40 \i_fifo_tx/U338  ( .A(\i_fifo_tx/mem[12][5] ), .B(
        \i_fifo_tx/mem[13][5] ), .C(\i_fifo_tx/mem[14][5] ), .D(
        \i_fifo_tx/mem[15][5] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n327 ) );
  IMUX40 \i_fifo_tx/U330  ( .A(\i_fifo_tx/mem[44][5] ), .B(
        \i_fifo_tx/mem[45][5] ), .C(\i_fifo_tx/mem[46][5] ), .D(
        \i_fifo_tx/mem[47][5] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n317 ) );
  IMUX40 \i_fifo_tx/U326  ( .A(\i_fifo_tx/mem[60][5] ), .B(
        \i_fifo_tx/mem[61][5] ), .C(\i_fifo_tx/mem[62][5] ), .D(
        \i_fifo_tx/mem[63][5] ), .S0(n315), .S1(n319), .Q(\i_fifo_tx/n312 ) );
  IMUX40 \i_fifo_tx/U350  ( .A(\i_fifo_tx/mem[28][6] ), .B(
        \i_fifo_tx/mem[29][6] ), .C(\i_fifo_tx/mem[30][6] ), .D(
        \i_fifo_tx/mem[31][6] ), .S0(n316), .S1(n318), .Q(\i_fifo_tx/n342 ) );
  IMUX40 \i_fifo_tx/U354  ( .A(\i_fifo_tx/mem[12][6] ), .B(
        \i_fifo_tx/mem[13][6] ), .C(\i_fifo_tx/mem[14][6] ), .D(
        \i_fifo_tx/mem[15][6] ), .S0(n132), .S1(n319), .Q(\i_fifo_tx/n347 ) );
  IMUX40 \i_fifo_tx/U346  ( .A(\i_fifo_tx/mem[44][6] ), .B(
        \i_fifo_tx/mem[45][6] ), .C(\i_fifo_tx/mem[46][6] ), .D(
        \i_fifo_tx/mem[47][6] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n337 ) );
  IMUX40 \i_fifo_tx/U342  ( .A(\i_fifo_tx/mem[60][6] ), .B(
        \i_fifo_tx/mem[61][6] ), .C(\i_fifo_tx/mem[62][6] ), .D(
        \i_fifo_tx/mem[63][6] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n332 ) );
  IMUX40 \i_fifo_tx/U366  ( .A(\i_fifo_tx/mem[28][7] ), .B(
        \i_fifo_tx/mem[29][7] ), .C(\i_fifo_tx/mem[30][7] ), .D(
        \i_fifo_tx/mem[31][7] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n362 ) );
  IMUX40 \i_fifo_tx/U373  ( .A(\i_fifo_tx/mem[0][7] ), .B(
        \i_fifo_tx/mem[1][7] ), .C(\i_fifo_tx/mem[2][7] ), .D(
        \i_fifo_tx/mem[3][7] ), .S0(n317), .S1(n318), .Q(\i_fifo_tx/n364 ) );
  IMUX40 \i_fifo_tx/U362  ( .A(\i_fifo_tx/mem[44][7] ), .B(
        \i_fifo_tx/mem[45][7] ), .C(\i_fifo_tx/mem[46][7] ), .D(
        \i_fifo_tx/mem[47][7] ), .S0(n315), .S1(n318), .Q(\i_fifo_tx/n357 ) );
  IMUX40 \i_fifo_tx/U358  ( .A(\i_fifo_tx/mem[60][7] ), .B(
        \i_fifo_tx/mem[61][7] ), .C(\i_fifo_tx/mem[62][7] ), .D(
        \i_fifo_tx/mem[63][7] ), .S0(n314), .S1(n319), .Q(\i_fifo_tx/n352 ) );
  IMUX40 \i_fifo_rx/U446  ( .A(\i_fifo_rx/mem[12][0] ), .B(
        \i_fifo_rx/mem[13][0] ), .C(\i_fifo_rx/mem[14][0] ), .D(
        \i_fifo_rx/mem[15][0] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n397 ) );
  IMUX40 \i_fifo_rx/U438  ( .A(\i_fifo_rx/mem[44][0] ), .B(
        \i_fifo_rx/mem[45][0] ), .C(\i_fifo_rx/mem[46][0] ), .D(
        \i_fifo_rx/mem[47][0] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n387 ) );
  IMUX40 \i_fifo_rx/U434  ( .A(\i_fifo_rx/mem[60][0] ), .B(
        \i_fifo_rx/mem[61][0] ), .C(\i_fifo_rx/mem[62][0] ), .D(
        \i_fifo_rx/mem[63][0] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n382 ) );
  IMUX40 \i_fifo_rx/U462  ( .A(\i_fifo_rx/mem[12][1] ), .B(
        \i_fifo_rx/mem[13][1] ), .C(\i_fifo_rx/mem[14][1] ), .D(
        \i_fifo_rx/mem[15][1] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n417 ) );
  IMUX40 \i_fifo_rx/U454  ( .A(\i_fifo_rx/mem[44][1] ), .B(
        \i_fifo_rx/mem[45][1] ), .C(\i_fifo_rx/mem[46][1] ), .D(
        \i_fifo_rx/mem[47][1] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n407 ) );
  IMUX40 \i_fifo_rx/U450  ( .A(\i_fifo_rx/mem[60][1] ), .B(
        \i_fifo_rx/mem[61][1] ), .C(\i_fifo_rx/mem[62][1] ), .D(
        \i_fifo_rx/mem[63][1] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n402 ) );
  IMUX40 \i_fifo_rx/U478  ( .A(\i_fifo_rx/mem[12][2] ), .B(
        \i_fifo_rx/mem[13][2] ), .C(\i_fifo_rx/mem[14][2] ), .D(
        \i_fifo_rx/mem[15][2] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n437 ) );
  IMUX40 \i_fifo_rx/U470  ( .A(\i_fifo_rx/mem[44][2] ), .B(
        \i_fifo_rx/mem[45][2] ), .C(\i_fifo_rx/mem[46][2] ), .D(
        \i_fifo_rx/mem[47][2] ), .S0(\i_fifo_rx/N39 ), .S1(n311), .Q(
        \i_fifo_rx/n427 ) );
  IMUX40 \i_fifo_rx/U466  ( .A(\i_fifo_rx/mem[60][2] ), .B(
        \i_fifo_rx/mem[61][2] ), .C(\i_fifo_rx/mem[62][2] ), .D(
        \i_fifo_rx/mem[63][2] ), .S0(\i_fifo_rx/N39 ), .S1(n311), .Q(
        \i_fifo_rx/n422 ) );
  IMUX40 \i_fifo_rx/U494  ( .A(\i_fifo_rx/mem[12][3] ), .B(
        \i_fifo_rx/mem[13][3] ), .C(\i_fifo_rx/mem[14][3] ), .D(
        \i_fifo_rx/mem[15][3] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n457 ) );
  IMUX40 \i_fifo_rx/U486  ( .A(\i_fifo_rx/mem[44][3] ), .B(
        \i_fifo_rx/mem[45][3] ), .C(\i_fifo_rx/mem[46][3] ), .D(
        \i_fifo_rx/mem[47][3] ), .S0(\i_fifo_rx/N39 ), .S1(n311), .Q(
        \i_fifo_rx/n447 ) );
  IMUX40 \i_fifo_rx/U482  ( .A(\i_fifo_rx/mem[60][3] ), .B(
        \i_fifo_rx/mem[61][3] ), .C(\i_fifo_rx/mem[62][3] ), .D(
        \i_fifo_rx/mem[63][3] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n442 ) );
  IMUX40 \i_fifo_rx/U510  ( .A(\i_fifo_rx/mem[12][4] ), .B(
        \i_fifo_rx/mem[13][4] ), .C(\i_fifo_rx/mem[14][4] ), .D(
        \i_fifo_rx/mem[15][4] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n477 ) );
  IMUX40 \i_fifo_rx/U502  ( .A(\i_fifo_rx/mem[44][4] ), .B(
        \i_fifo_rx/mem[45][4] ), .C(\i_fifo_rx/mem[46][4] ), .D(
        \i_fifo_rx/mem[47][4] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n467 ) );
  IMUX40 \i_fifo_rx/U498  ( .A(\i_fifo_rx/mem[60][4] ), .B(
        \i_fifo_rx/mem[61][4] ), .C(\i_fifo_rx/mem[62][4] ), .D(
        \i_fifo_rx/mem[63][4] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n462 ) );
  IMUX40 \i_fifo_rx/U526  ( .A(\i_fifo_rx/mem[12][5] ), .B(
        \i_fifo_rx/mem[13][5] ), .C(\i_fifo_rx/mem[14][5] ), .D(
        \i_fifo_rx/mem[15][5] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n497 ) );
  IMUX40 \i_fifo_rx/U518  ( .A(\i_fifo_rx/mem[44][5] ), .B(
        \i_fifo_rx/mem[45][5] ), .C(\i_fifo_rx/mem[46][5] ), .D(
        \i_fifo_rx/mem[47][5] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n487 ) );
  IMUX40 \i_fifo_rx/U514  ( .A(\i_fifo_rx/mem[60][5] ), .B(
        \i_fifo_rx/mem[61][5] ), .C(\i_fifo_rx/mem[62][5] ), .D(
        \i_fifo_rx/mem[63][5] ), .S0(\i_fifo_rx/N39 ), .S1(n311), .Q(
        \i_fifo_rx/n482 ) );
  IMUX40 \i_fifo_rx/U542  ( .A(\i_fifo_rx/mem[12][6] ), .B(
        \i_fifo_rx/mem[13][6] ), .C(\i_fifo_rx/mem[14][6] ), .D(
        \i_fifo_rx/mem[15][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n517 ) );
  IMUX40 \i_fifo_rx/U534  ( .A(\i_fifo_rx/mem[44][6] ), .B(
        \i_fifo_rx/mem[45][6] ), .C(\i_fifo_rx/mem[46][6] ), .D(
        \i_fifo_rx/mem[47][6] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n507 ) );
  IMUX40 \i_fifo_rx/U530  ( .A(\i_fifo_rx/mem[60][6] ), .B(
        \i_fifo_rx/mem[61][6] ), .C(\i_fifo_rx/mem[62][6] ), .D(
        \i_fifo_rx/mem[63][6] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n502 ) );
  IMUX40 \i_fifo_rx/U558  ( .A(\i_fifo_rx/mem[12][7] ), .B(
        \i_fifo_rx/mem[13][7] ), .C(\i_fifo_rx/mem[14][7] ), .D(
        \i_fifo_rx/mem[15][7] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n537 ) );
  IMUX40 \i_fifo_rx/U550  ( .A(\i_fifo_rx/mem[44][7] ), .B(
        \i_fifo_rx/mem[45][7] ), .C(\i_fifo_rx/mem[46][7] ), .D(
        \i_fifo_rx/mem[47][7] ), .S0(n306), .S1(n311), .Q(\i_fifo_rx/n527 ) );
  IMUX40 \i_fifo_rx/U546  ( .A(\i_fifo_rx/mem[60][7] ), .B(
        \i_fifo_rx/mem[61][7] ), .C(\i_fifo_rx/mem[62][7] ), .D(
        \i_fifo_rx/mem[63][7] ), .S0(n307), .S1(n311), .Q(\i_fifo_rx/n522 ) );
  IMUX40 \i_fifo_rx/U278  ( .A(\i_fifo_rx/mem[12][0] ), .B(
        \i_fifo_rx/mem[13][0] ), .C(\i_fifo_rx/mem[14][0] ), .D(
        \i_fifo_rx/mem[15][0] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n237 ) );
  IMUX40 \i_fifo_rx/U270  ( .A(\i_fifo_rx/mem[44][0] ), .B(
        \i_fifo_rx/mem[45][0] ), .C(\i_fifo_rx/mem[46][0] ), .D(
        \i_fifo_rx/mem[47][0] ), .S0(n302), .S1(n303), .Q(\i_fifo_rx/n227 ) );
  IMUX40 \i_fifo_rx/U266  ( .A(\i_fifo_rx/mem[60][0] ), .B(
        \i_fifo_rx/mem[61][0] ), .C(\i_fifo_rx/mem[62][0] ), .D(
        \i_fifo_rx/mem[63][0] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n222 ) );
  IMUX40 \i_fifo_rx/U294  ( .A(\i_fifo_rx/mem[12][1] ), .B(
        \i_fifo_rx/mem[13][1] ), .C(\i_fifo_rx/mem[14][1] ), .D(
        \i_fifo_rx/mem[15][1] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n257 ) );
  IMUX40 \i_fifo_rx/U286  ( .A(\i_fifo_rx/mem[44][1] ), .B(
        \i_fifo_rx/mem[45][1] ), .C(\i_fifo_rx/mem[46][1] ), .D(
        \i_fifo_rx/mem[47][1] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n247 ) );
  IMUX40 \i_fifo_rx/U282  ( .A(\i_fifo_rx/mem[60][1] ), .B(
        \i_fifo_rx/mem[61][1] ), .C(\i_fifo_rx/mem[62][1] ), .D(
        \i_fifo_rx/mem[63][1] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n242 ) );
  IMUX40 \i_fifo_rx/U310  ( .A(\i_fifo_rx/mem[12][2] ), .B(
        \i_fifo_rx/mem[13][2] ), .C(\i_fifo_rx/mem[14][2] ), .D(
        \i_fifo_rx/mem[15][2] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n277 ) );
  IMUX40 \i_fifo_rx/U302  ( .A(\i_fifo_rx/mem[44][2] ), .B(
        \i_fifo_rx/mem[45][2] ), .C(\i_fifo_rx/mem[46][2] ), .D(
        \i_fifo_rx/mem[47][2] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n267 ) );
  IMUX40 \i_fifo_rx/U298  ( .A(\i_fifo_rx/mem[60][2] ), .B(
        \i_fifo_rx/mem[61][2] ), .C(\i_fifo_rx/mem[62][2] ), .D(
        \i_fifo_rx/mem[63][2] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n262 ) );
  IMUX40 \i_fifo_rx/U326  ( .A(\i_fifo_rx/mem[12][3] ), .B(
        \i_fifo_rx/mem[13][3] ), .C(\i_fifo_rx/mem[14][3] ), .D(
        \i_fifo_rx/mem[15][3] ), .S0(n299), .S1(n305), .Q(\i_fifo_rx/n297 ) );
  IMUX40 \i_fifo_rx/U318  ( .A(\i_fifo_rx/mem[44][3] ), .B(
        \i_fifo_rx/mem[45][3] ), .C(\i_fifo_rx/mem[46][3] ), .D(
        \i_fifo_rx/mem[47][3] ), .S0(n134), .S1(n305), .Q(\i_fifo_rx/n287 ) );
  IMUX40 \i_fifo_rx/U314  ( .A(\i_fifo_rx/mem[60][3] ), .B(
        \i_fifo_rx/mem[61][3] ), .C(\i_fifo_rx/mem[62][3] ), .D(
        \i_fifo_rx/mem[63][3] ), .S0(n134), .S1(n305), .Q(\i_fifo_rx/n282 ) );
  IMUX40 \i_fifo_rx/U342  ( .A(\i_fifo_rx/mem[12][4] ), .B(
        \i_fifo_rx/mem[13][4] ), .C(\i_fifo_rx/mem[14][4] ), .D(
        \i_fifo_rx/mem[15][4] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n317 ) );
  IMUX40 \i_fifo_rx/U334  ( .A(\i_fifo_rx/mem[44][4] ), .B(
        \i_fifo_rx/mem[45][4] ), .C(\i_fifo_rx/mem[46][4] ), .D(
        \i_fifo_rx/mem[47][4] ), .S0(n134), .S1(n305), .Q(\i_fifo_rx/n307 ) );
  IMUX40 \i_fifo_rx/U330  ( .A(\i_fifo_rx/mem[60][4] ), .B(
        \i_fifo_rx/mem[61][4] ), .C(\i_fifo_rx/mem[62][4] ), .D(
        \i_fifo_rx/mem[63][4] ), .S0(n300), .S1(n305), .Q(\i_fifo_rx/n302 ) );
  IMUX40 \i_fifo_rx/U358  ( .A(\i_fifo_rx/mem[12][5] ), .B(
        \i_fifo_rx/mem[13][5] ), .C(\i_fifo_rx/mem[14][5] ), .D(
        \i_fifo_rx/mem[15][5] ), .S0(n300), .S1(n86), .Q(\i_fifo_rx/n337 ) );
  IMUX40 \i_fifo_rx/U350  ( .A(\i_fifo_rx/mem[44][5] ), .B(
        \i_fifo_rx/mem[45][5] ), .C(\i_fifo_rx/mem[46][5] ), .D(
        \i_fifo_rx/mem[47][5] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n327 ) );
  IMUX40 \i_fifo_rx/U346  ( .A(\i_fifo_rx/mem[60][5] ), .B(
        \i_fifo_rx/mem[61][5] ), .C(\i_fifo_rx/mem[62][5] ), .D(
        \i_fifo_rx/mem[63][5] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n322 ) );
  IMUX40 \i_fifo_rx/U374  ( .A(\i_fifo_rx/mem[12][6] ), .B(
        \i_fifo_rx/mem[13][6] ), .C(\i_fifo_rx/mem[14][6] ), .D(
        \i_fifo_rx/mem[15][6] ), .S0(n134), .S1(n303), .Q(\i_fifo_rx/n357 ) );
  IMUX40 \i_fifo_rx/U366  ( .A(\i_fifo_rx/mem[44][6] ), .B(
        \i_fifo_rx/mem[45][6] ), .C(\i_fifo_rx/mem[46][6] ), .D(
        \i_fifo_rx/mem[47][6] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n347 ) );
  IMUX40 \i_fifo_rx/U362  ( .A(\i_fifo_rx/mem[60][6] ), .B(
        \i_fifo_rx/mem[61][6] ), .C(\i_fifo_rx/mem[62][6] ), .D(
        \i_fifo_rx/mem[63][6] ), .S0(n300), .S1(n303), .Q(\i_fifo_rx/n342 ) );
  IMUX40 \i_fifo_rx/U393  ( .A(\i_fifo_rx/mem[0][7] ), .B(
        \i_fifo_rx/mem[1][7] ), .C(\i_fifo_rx/mem[2][7] ), .D(
        \i_fifo_rx/mem[3][7] ), .S0(n302), .S1(n305), .Q(\i_fifo_rx/n374 ) );
  IMUX40 \i_fifo_rx/U382  ( .A(\i_fifo_rx/mem[44][7] ), .B(
        \i_fifo_rx/mem[45][7] ), .C(\i_fifo_rx/mem[46][7] ), .D(
        \i_fifo_rx/mem[47][7] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n367 ) );
  IMUX40 \i_fifo_rx/U378  ( .A(\i_fifo_rx/mem[60][7] ), .B(
        \i_fifo_rx/mem[61][7] ), .C(\i_fifo_rx/mem[62][7] ), .D(
        \i_fifo_rx/mem[63][7] ), .S0(n299), .S1(n303), .Q(\i_fifo_rx/n362 ) );
  MUX41 \i_fifo_tx/U383  ( .A(\i_fifo_tx/n403 ), .B(\i_fifo_tx/n393 ), .C(
        \i_fifo_tx/n398 ), .D(\i_fifo_tx/n388 ), .S0(\i_fifo_tx/N35 ), .S1(
        \i_fifo_tx/N34 ), .Q(\i_fifo_tx/N142 ) );
  MUX41 \i_fifo_tx/U378  ( .A(\i_fifo_tx/n383 ), .B(\i_fifo_tx/n373 ), .C(
        \i_fifo_tx/n378 ), .D(\i_fifo_tx/n368 ), .S0(\i_fifo_tx/N35 ), .S1(
        \i_fifo_tx/N34 ), .Q(\i_fifo_tx/N143 ) );
  MUX41 \i_fifo_tx/U388  ( .A(\i_fifo_tx/n423 ), .B(\i_fifo_tx/n413 ), .C(
        \i_fifo_tx/n418 ), .D(\i_fifo_tx/n408 ), .S0(\i_fifo_tx/N35 ), .S1(
        \i_fifo_tx/N34 ), .Q(\i_fifo_tx/N141 ) );
  IMUX40 \i_fifo_tx/U544  ( .A(\i_fifo_tx/N143 ), .B(\i_fifo_tx/N142 ), .C(
        \i_fifo_tx/N141 ), .D(\i_fifo_tx/N140 ), .S0(\i_fifo_tx/N36 ), .S1(
        \i_fifo_tx/N37 ), .Q(\i_fifo_tx/n528 ) );
  MUX41 \i_fifo_tx/U403  ( .A(\i_fifo_tx/n483 ), .B(\i_fifo_tx/n473 ), .C(
        \i_fifo_tx/n478 ), .D(\i_fifo_tx/n468 ), .S0(\i_fifo_tx/N35 ), .S1(
        \i_fifo_tx/N34 ), .Q(\i_fifo_tx/N138 ) );
  MUX41 \i_fifo_tx/U398  ( .A(\i_fifo_tx/n463 ), .B(\i_fifo_tx/n453 ), .C(
        \i_fifo_tx/n458 ), .D(\i_fifo_tx/n448 ), .S0(\i_fifo_tx/N35 ), .S1(
        \i_fifo_tx/N34 ), .Q(\i_fifo_tx/N139 ) );
  MUX41 \i_fifo_tx/U408  ( .A(\i_fifo_tx/n503 ), .B(\i_fifo_tx/n493 ), .C(
        \i_fifo_tx/n498 ), .D(\i_fifo_tx/n488 ), .S0(\i_fifo_tx/N35 ), .S1(
        \i_fifo_tx/N34 ), .Q(\i_fifo_tx/N137 ) );
  IMUX40 \i_fifo_tx/U543  ( .A(\i_fifo_tx/N139 ), .B(\i_fifo_tx/N138 ), .C(
        \i_fifo_tx/N137 ), .D(\i_fifo_tx/N136 ), .S0(\i_fifo_tx/N36 ), .S1(
        \i_fifo_tx/N37 ), .Q(\i_fifo_tx/n529 ) );
  IMUX40 \i_fifo_tx/U390  ( .A(\i_fifo_tx/n434 ), .B(\i_fifo_tx/n435 ), .C(
        \i_fifo_tx/n436 ), .D(\i_fifo_tx/n437 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n433 ) );
  IMUX40 \i_fifo_tx/U392  ( .A(\i_fifo_tx/n444 ), .B(\i_fifo_tx/n445 ), .C(
        \i_fifo_tx/n446 ), .D(\i_fifo_tx/n447 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n443 ) );
  IMUX40 \i_fifo_tx/U391  ( .A(\i_fifo_tx/n439 ), .B(\i_fifo_tx/n440 ), .C(
        \i_fifo_tx/n441 ), .D(\i_fifo_tx/n442 ), .S0(\i_fifo_tx/N33 ), .S1(
        n1941), .Q(\i_fifo_tx/n438 ) );
  MUX41 \i_fifo_tx/U393  ( .A(\i_fifo_tx/n443 ), .B(\i_fifo_tx/n433 ), .C(
        \i_fifo_tx/n438 ), .D(\i_fifo_tx/n428 ), .S0(\i_fifo_tx/N35 ), .S1(
        \i_fifo_tx/N34 ), .Q(\i_fifo_tx/N140 ) );
  IMUX40 \i_fifo_tx/U455  ( .A(\i_fifo_tx/mem[24][2] ), .B(
        \i_fifo_tx/mem[25][2] ), .C(\i_fifo_tx/mem[26][2] ), .D(
        \i_fifo_tx/mem[27][2] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n420 ) );
  IMUX40 \i_fifo_tx/U457  ( .A(\i_fifo_tx/mem[16][2] ), .B(
        \i_fifo_tx/mem[17][2] ), .C(\i_fifo_tx/mem[18][2] ), .D(
        \i_fifo_tx/mem[19][2] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n419 ) );
  IMUX40 \i_fifo_tx/U456  ( .A(\i_fifo_tx/mem[20][2] ), .B(
        \i_fifo_tx/mem[21][2] ), .C(\i_fifo_tx/mem[22][2] ), .D(
        \i_fifo_tx/mem[23][2] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n421 ) );
  IMUX40 \i_fifo_tx/U386  ( .A(\i_fifo_tx/n419 ), .B(\i_fifo_tx/n420 ), .C(
        \i_fifo_tx/n421 ), .D(\i_fifo_tx/n422 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n418 ) );
  IMUX40 \i_fifo_tx/U459  ( .A(\i_fifo_tx/mem[8][2] ), .B(
        \i_fifo_tx/mem[9][2] ), .C(\i_fifo_tx/mem[10][2] ), .D(
        \i_fifo_tx/mem[11][2] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n425 ) );
  IMUX40 \i_fifo_tx/U461  ( .A(\i_fifo_tx/mem[0][2] ), .B(
        \i_fifo_tx/mem[1][2] ), .C(\i_fifo_tx/mem[2][2] ), .D(
        \i_fifo_tx/mem[3][2] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n424 ) );
  IMUX40 \i_fifo_tx/U460  ( .A(\i_fifo_tx/mem[4][2] ), .B(
        \i_fifo_tx/mem[5][2] ), .C(\i_fifo_tx/mem[6][2] ), .D(
        \i_fifo_tx/mem[7][2] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n426 ) );
  IMUX40 \i_fifo_tx/U387  ( .A(\i_fifo_tx/n424 ), .B(\i_fifo_tx/n425 ), .C(
        \i_fifo_tx/n426 ), .D(\i_fifo_tx/n427 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n423 ) );
  IMUX40 \i_fifo_tx/U451  ( .A(\i_fifo_tx/mem[40][2] ), .B(
        \i_fifo_tx/mem[41][2] ), .C(\i_fifo_tx/mem[42][2] ), .D(
        \i_fifo_tx/mem[43][2] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n415 ) );
  IMUX40 \i_fifo_tx/U453  ( .A(\i_fifo_tx/mem[32][2] ), .B(
        \i_fifo_tx/mem[33][2] ), .C(\i_fifo_tx/mem[34][2] ), .D(
        \i_fifo_tx/mem[35][2] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n414 ) );
  IMUX40 \i_fifo_tx/U452  ( .A(\i_fifo_tx/mem[36][2] ), .B(
        \i_fifo_tx/mem[37][2] ), .C(\i_fifo_tx/mem[38][2] ), .D(
        \i_fifo_tx/mem[39][2] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n416 ) );
  IMUX40 \i_fifo_tx/U385  ( .A(\i_fifo_tx/n414 ), .B(\i_fifo_tx/n415 ), .C(
        \i_fifo_tx/n416 ), .D(\i_fifo_tx/n417 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n413 ) );
  IMUX40 \i_fifo_tx/U447  ( .A(\i_fifo_tx/mem[56][2] ), .B(
        \i_fifo_tx/mem[57][2] ), .C(\i_fifo_tx/mem[58][2] ), .D(
        \i_fifo_tx/mem[59][2] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n410 ) );
  IMUX40 \i_fifo_tx/U449  ( .A(\i_fifo_tx/mem[48][2] ), .B(
        \i_fifo_tx/mem[49][2] ), .C(\i_fifo_tx/mem[50][2] ), .D(
        \i_fifo_tx/mem[51][2] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n409 ) );
  IMUX40 \i_fifo_tx/U448  ( .A(\i_fifo_tx/mem[52][2] ), .B(
        \i_fifo_tx/mem[53][2] ), .C(\i_fifo_tx/mem[54][2] ), .D(
        \i_fifo_tx/mem[55][2] ), .S0(n324), .S1(\i_fifo_tx/N31 ), .Q(
        \i_fifo_tx/n411 ) );
  IMUX40 \i_fifo_tx/U384  ( .A(\i_fifo_tx/n409 ), .B(\i_fifo_tx/n410 ), .C(
        \i_fifo_tx/n411 ), .D(\i_fifo_tx/n412 ), .S0(n270), .S1(
        \i_fifo_tx/N32 ), .Q(\i_fifo_tx/n408 ) );
  IMUX40 \i_fifo_tx/U423  ( .A(\i_fifo_tx/mem[24][0] ), .B(
        \i_fifo_tx/mem[25][0] ), .C(\i_fifo_tx/mem[26][0] ), .D(
        \i_fifo_tx/mem[27][0] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n380 ) );
  IMUX40 \i_fifo_tx/U425  ( .A(\i_fifo_tx/mem[16][0] ), .B(
        \i_fifo_tx/mem[17][0] ), .C(\i_fifo_tx/mem[18][0] ), .D(
        \i_fifo_tx/mem[19][0] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n379 ) );
  IMUX40 \i_fifo_tx/U424  ( .A(\i_fifo_tx/mem[20][0] ), .B(
        \i_fifo_tx/mem[21][0] ), .C(\i_fifo_tx/mem[22][0] ), .D(
        \i_fifo_tx/mem[23][0] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n381 ) );
  IMUX40 \i_fifo_tx/U376  ( .A(\i_fifo_tx/n379 ), .B(\i_fifo_tx/n380 ), .C(
        \i_fifo_tx/n381 ), .D(\i_fifo_tx/n382 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n378 ) );
  IMUX40 \i_fifo_tx/U427  ( .A(\i_fifo_tx/mem[8][0] ), .B(
        \i_fifo_tx/mem[9][0] ), .C(\i_fifo_tx/mem[10][0] ), .D(
        \i_fifo_tx/mem[11][0] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n385 ) );
  IMUX40 \i_fifo_tx/U429  ( .A(\i_fifo_tx/mem[0][0] ), .B(
        \i_fifo_tx/mem[1][0] ), .C(\i_fifo_tx/mem[2][0] ), .D(
        \i_fifo_tx/mem[3][0] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n384 ) );
  IMUX40 \i_fifo_tx/U428  ( .A(\i_fifo_tx/mem[4][0] ), .B(
        \i_fifo_tx/mem[5][0] ), .C(\i_fifo_tx/mem[6][0] ), .D(
        \i_fifo_tx/mem[7][0] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n386 ) );
  IMUX40 \i_fifo_tx/U377  ( .A(\i_fifo_tx/n384 ), .B(\i_fifo_tx/n385 ), .C(
        \i_fifo_tx/n386 ), .D(\i_fifo_tx/n387 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n383 ) );
  IMUX40 \i_fifo_tx/U419  ( .A(\i_fifo_tx/mem[40][0] ), .B(
        \i_fifo_tx/mem[41][0] ), .C(\i_fifo_tx/mem[42][0] ), .D(
        \i_fifo_tx/mem[43][0] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n375 ) );
  IMUX40 \i_fifo_tx/U421  ( .A(\i_fifo_tx/mem[32][0] ), .B(
        \i_fifo_tx/mem[33][0] ), .C(\i_fifo_tx/mem[34][0] ), .D(
        \i_fifo_tx/mem[35][0] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n374 ) );
  IMUX40 \i_fifo_tx/U420  ( .A(\i_fifo_tx/mem[36][0] ), .B(
        \i_fifo_tx/mem[37][0] ), .C(\i_fifo_tx/mem[38][0] ), .D(
        \i_fifo_tx/mem[39][0] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n376 ) );
  IMUX40 \i_fifo_tx/U375  ( .A(\i_fifo_tx/n374 ), .B(\i_fifo_tx/n375 ), .C(
        \i_fifo_tx/n376 ), .D(\i_fifo_tx/n377 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n373 ) );
  IMUX40 \i_fifo_tx/U415  ( .A(\i_fifo_tx/mem[56][0] ), .B(
        \i_fifo_tx/mem[57][0] ), .C(\i_fifo_tx/mem[58][0] ), .D(
        \i_fifo_tx/mem[59][0] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n370 ) );
  IMUX40 \i_fifo_tx/U417  ( .A(\i_fifo_tx/mem[48][0] ), .B(
        \i_fifo_tx/mem[49][0] ), .C(\i_fifo_tx/mem[50][0] ), .D(
        \i_fifo_tx/mem[51][0] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n369 ) );
  IMUX40 \i_fifo_tx/U416  ( .A(\i_fifo_tx/mem[52][0] ), .B(
        \i_fifo_tx/mem[53][0] ), .C(\i_fifo_tx/mem[54][0] ), .D(
        \i_fifo_tx/mem[55][0] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n371 ) );
  IMUX40 \i_fifo_tx/U374  ( .A(\i_fifo_tx/n369 ), .B(\i_fifo_tx/n370 ), .C(
        \i_fifo_tx/n371 ), .D(\i_fifo_tx/n372 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n368 ) );
  IMUX40 \i_fifo_tx/U439  ( .A(\i_fifo_tx/mem[24][1] ), .B(
        \i_fifo_tx/mem[25][1] ), .C(\i_fifo_tx/mem[26][1] ), .D(
        \i_fifo_tx/mem[27][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n400 ) );
  IMUX40 \i_fifo_tx/U441  ( .A(\i_fifo_tx/mem[16][1] ), .B(
        \i_fifo_tx/mem[17][1] ), .C(\i_fifo_tx/mem[18][1] ), .D(
        \i_fifo_tx/mem[19][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n399 ) );
  IMUX40 \i_fifo_tx/U440  ( .A(\i_fifo_tx/mem[20][1] ), .B(
        \i_fifo_tx/mem[21][1] ), .C(\i_fifo_tx/mem[22][1] ), .D(
        \i_fifo_tx/mem[23][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n401 ) );
  IMUX40 \i_fifo_tx/U381  ( .A(\i_fifo_tx/n399 ), .B(\i_fifo_tx/n400 ), .C(
        \i_fifo_tx/n401 ), .D(\i_fifo_tx/n402 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n398 ) );
  IMUX40 \i_fifo_tx/U443  ( .A(\i_fifo_tx/mem[8][1] ), .B(
        \i_fifo_tx/mem[9][1] ), .C(\i_fifo_tx/mem[10][1] ), .D(
        \i_fifo_tx/mem[11][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n405 ) );
  IMUX40 \i_fifo_tx/U445  ( .A(\i_fifo_tx/mem[0][1] ), .B(
        \i_fifo_tx/mem[1][1] ), .C(\i_fifo_tx/mem[2][1] ), .D(
        \i_fifo_tx/mem[3][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n404 ) );
  IMUX40 \i_fifo_tx/U444  ( .A(\i_fifo_tx/mem[4][1] ), .B(
        \i_fifo_tx/mem[5][1] ), .C(\i_fifo_tx/mem[6][1] ), .D(
        \i_fifo_tx/mem[7][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n406 ) );
  IMUX40 \i_fifo_tx/U382  ( .A(\i_fifo_tx/n404 ), .B(\i_fifo_tx/n405 ), .C(
        \i_fifo_tx/n406 ), .D(\i_fifo_tx/n407 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n403 ) );
  IMUX40 \i_fifo_tx/U435  ( .A(\i_fifo_tx/mem[40][1] ), .B(
        \i_fifo_tx/mem[41][1] ), .C(\i_fifo_tx/mem[42][1] ), .D(
        \i_fifo_tx/mem[43][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n395 ) );
  IMUX40 \i_fifo_tx/U437  ( .A(\i_fifo_tx/mem[32][1] ), .B(
        \i_fifo_tx/mem[33][1] ), .C(\i_fifo_tx/mem[34][1] ), .D(
        \i_fifo_tx/mem[35][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n394 ) );
  IMUX40 \i_fifo_tx/U436  ( .A(\i_fifo_tx/mem[36][1] ), .B(
        \i_fifo_tx/mem[37][1] ), .C(\i_fifo_tx/mem[38][1] ), .D(
        \i_fifo_tx/mem[39][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n396 ) );
  IMUX40 \i_fifo_tx/U380  ( .A(\i_fifo_tx/n394 ), .B(\i_fifo_tx/n395 ), .C(
        \i_fifo_tx/n396 ), .D(\i_fifo_tx/n397 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n393 ) );
  IMUX40 \i_fifo_tx/U431  ( .A(\i_fifo_tx/mem[56][1] ), .B(
        \i_fifo_tx/mem[57][1] ), .C(\i_fifo_tx/mem[58][1] ), .D(
        \i_fifo_tx/mem[59][1] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n390 ) );
  IMUX40 \i_fifo_tx/U433  ( .A(\i_fifo_tx/mem[48][1] ), .B(
        \i_fifo_tx/mem[49][1] ), .C(\i_fifo_tx/mem[50][1] ), .D(
        \i_fifo_tx/mem[51][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n389 ) );
  IMUX40 \i_fifo_tx/U432  ( .A(\i_fifo_tx/mem[52][1] ), .B(
        \i_fifo_tx/mem[53][1] ), .C(\i_fifo_tx/mem[54][1] ), .D(
        \i_fifo_tx/mem[55][1] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n391 ) );
  IMUX40 \i_fifo_tx/U379  ( .A(\i_fifo_tx/n389 ), .B(\i_fifo_tx/n390 ), .C(
        \i_fifo_tx/n391 ), .D(\i_fifo_tx/n392 ), .S0(\i_fifo_tx/N33 ), .S1(
        \i_fifo_tx/N32 ), .Q(\i_fifo_tx/n388 ) );
  IMUX40 \i_fifo_tx/U410  ( .A(\i_fifo_tx/n514 ), .B(\i_fifo_tx/n515 ), .C(
        \i_fifo_tx/n516 ), .D(\i_fifo_tx/n517 ), .S0(\i_fifo_tx/N33 ), .S1(
        \i_fifo_tx/N32 ), .Q(\i_fifo_tx/n513 ) );
  IMUX40 \i_fifo_tx/U412  ( .A(\i_fifo_tx/n524 ), .B(\i_fifo_tx/n525 ), .C(
        \i_fifo_tx/n526 ), .D(\i_fifo_tx/n527 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n523 ) );
  IMUX40 \i_fifo_tx/U411  ( .A(\i_fifo_tx/n519 ), .B(\i_fifo_tx/n520 ), .C(
        \i_fifo_tx/n521 ), .D(\i_fifo_tx/n522 ), .S0(\i_fifo_tx/N33 ), .S1(
        \i_fifo_tx/N32 ), .Q(\i_fifo_tx/n518 ) );
  MUX41 \i_fifo_tx/U413  ( .A(\i_fifo_tx/n523 ), .B(\i_fifo_tx/n513 ), .C(
        \i_fifo_tx/n518 ), .D(\i_fifo_tx/n508 ), .S0(\i_fifo_tx/N35 ), .S1(
        \i_fifo_tx/N34 ), .Q(\i_fifo_tx/N136 ) );
  IMUX40 \i_fifo_tx/U519  ( .A(\i_fifo_tx/mem[24][6] ), .B(
        \i_fifo_tx/mem[25][6] ), .C(\i_fifo_tx/mem[26][6] ), .D(
        \i_fifo_tx/mem[27][6] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n500 ) );
  IMUX40 \i_fifo_tx/U521  ( .A(\i_fifo_tx/mem[16][6] ), .B(
        \i_fifo_tx/mem[17][6] ), .C(\i_fifo_tx/mem[18][6] ), .D(
        \i_fifo_tx/mem[19][6] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n499 ) );
  IMUX40 \i_fifo_tx/U520  ( .A(\i_fifo_tx/mem[20][6] ), .B(
        \i_fifo_tx/mem[21][6] ), .C(\i_fifo_tx/mem[22][6] ), .D(
        \i_fifo_tx/mem[23][6] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n501 ) );
  IMUX40 \i_fifo_tx/U406  ( .A(\i_fifo_tx/n499 ), .B(\i_fifo_tx/n500 ), .C(
        \i_fifo_tx/n501 ), .D(\i_fifo_tx/n502 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n498 ) );
  IMUX40 \i_fifo_tx/U523  ( .A(\i_fifo_tx/mem[8][6] ), .B(
        \i_fifo_tx/mem[9][6] ), .C(\i_fifo_tx/mem[10][6] ), .D(
        \i_fifo_tx/mem[11][6] ), .S0(n321), .S1(\i_fifo_tx/N31 ), .Q(
        \i_fifo_tx/n505 ) );
  IMUX40 \i_fifo_tx/U525  ( .A(\i_fifo_tx/mem[0][6] ), .B(
        \i_fifo_tx/mem[1][6] ), .C(\i_fifo_tx/mem[2][6] ), .D(
        \i_fifo_tx/mem[3][6] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n504 ) );
  IMUX40 \i_fifo_tx/U524  ( .A(\i_fifo_tx/mem[4][6] ), .B(
        \i_fifo_tx/mem[5][6] ), .C(\i_fifo_tx/mem[6][6] ), .D(
        \i_fifo_tx/mem[7][6] ), .S0(n324), .S1(\i_fifo_tx/N31 ), .Q(
        \i_fifo_tx/n506 ) );
  IMUX40 \i_fifo_tx/U407  ( .A(\i_fifo_tx/n504 ), .B(\i_fifo_tx/n505 ), .C(
        \i_fifo_tx/n506 ), .D(\i_fifo_tx/n507 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n503 ) );
  IMUX40 \i_fifo_tx/U515  ( .A(\i_fifo_tx/mem[40][6] ), .B(
        \i_fifo_tx/mem[41][6] ), .C(\i_fifo_tx/mem[42][6] ), .D(
        \i_fifo_tx/mem[43][6] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n495 ) );
  IMUX40 \i_fifo_tx/U517  ( .A(\i_fifo_tx/mem[32][6] ), .B(
        \i_fifo_tx/mem[33][6] ), .C(\i_fifo_tx/mem[34][6] ), .D(
        \i_fifo_tx/mem[35][6] ), .S0(n324), .S1(\i_fifo_tx/N31 ), .Q(
        \i_fifo_tx/n494 ) );
  IMUX40 \i_fifo_tx/U516  ( .A(\i_fifo_tx/mem[36][6] ), .B(
        \i_fifo_tx/mem[37][6] ), .C(\i_fifo_tx/mem[38][6] ), .D(
        \i_fifo_tx/mem[39][6] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n496 ) );
  IMUX40 \i_fifo_tx/U405  ( .A(\i_fifo_tx/n494 ), .B(\i_fifo_tx/n495 ), .C(
        \i_fifo_tx/n496 ), .D(\i_fifo_tx/n497 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n493 ) );
  IMUX40 \i_fifo_tx/U511  ( .A(\i_fifo_tx/mem[56][6] ), .B(
        \i_fifo_tx/mem[57][6] ), .C(\i_fifo_tx/mem[58][6] ), .D(
        \i_fifo_tx/mem[59][6] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n490 ) );
  IMUX40 \i_fifo_tx/U513  ( .A(\i_fifo_tx/mem[48][6] ), .B(
        \i_fifo_tx/mem[49][6] ), .C(\i_fifo_tx/mem[50][6] ), .D(
        \i_fifo_tx/mem[51][6] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n489 ) );
  IMUX40 \i_fifo_tx/U512  ( .A(\i_fifo_tx/mem[52][6] ), .B(
        \i_fifo_tx/mem[53][6] ), .C(\i_fifo_tx/mem[54][6] ), .D(
        \i_fifo_tx/mem[55][6] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n491 ) );
  IMUX40 \i_fifo_tx/U404  ( .A(\i_fifo_tx/n489 ), .B(\i_fifo_tx/n490 ), .C(
        \i_fifo_tx/n491 ), .D(\i_fifo_tx/n492 ), .S0(\i_fifo_tx/N33 ), .S1(
        \i_fifo_tx/N32 ), .Q(\i_fifo_tx/n488 ) );
  IMUX40 \i_fifo_tx/U487  ( .A(\i_fifo_tx/mem[24][4] ), .B(
        \i_fifo_tx/mem[25][4] ), .C(\i_fifo_tx/mem[26][4] ), .D(
        \i_fifo_tx/mem[27][4] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n460 ) );
  IMUX40 \i_fifo_tx/U489  ( .A(\i_fifo_tx/mem[16][4] ), .B(
        \i_fifo_tx/mem[17][4] ), .C(\i_fifo_tx/mem[18][4] ), .D(
        \i_fifo_tx/mem[19][4] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n459 ) );
  IMUX40 \i_fifo_tx/U488  ( .A(\i_fifo_tx/mem[20][4] ), .B(
        \i_fifo_tx/mem[21][4] ), .C(\i_fifo_tx/mem[22][4] ), .D(
        \i_fifo_tx/mem[23][4] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n461 ) );
  IMUX40 \i_fifo_tx/U396  ( .A(\i_fifo_tx/n459 ), .B(\i_fifo_tx/n460 ), .C(
        \i_fifo_tx/n461 ), .D(\i_fifo_tx/n462 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n458 ) );
  IMUX40 \i_fifo_tx/U491  ( .A(\i_fifo_tx/mem[8][4] ), .B(
        \i_fifo_tx/mem[9][4] ), .C(\i_fifo_tx/mem[10][4] ), .D(
        \i_fifo_tx/mem[11][4] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n465 ) );
  IMUX40 \i_fifo_tx/U493  ( .A(\i_fifo_tx/mem[0][4] ), .B(
        \i_fifo_tx/mem[1][4] ), .C(\i_fifo_tx/mem[2][4] ), .D(
        \i_fifo_tx/mem[3][4] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n464 ) );
  IMUX40 \i_fifo_tx/U492  ( .A(\i_fifo_tx/mem[4][4] ), .B(
        \i_fifo_tx/mem[5][4] ), .C(\i_fifo_tx/mem[6][4] ), .D(
        \i_fifo_tx/mem[7][4] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n466 ) );
  IMUX40 \i_fifo_tx/U397  ( .A(\i_fifo_tx/n464 ), .B(\i_fifo_tx/n465 ), .C(
        \i_fifo_tx/n466 ), .D(\i_fifo_tx/n467 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n463 ) );
  IMUX40 \i_fifo_tx/U483  ( .A(\i_fifo_tx/mem[40][4] ), .B(
        \i_fifo_tx/mem[41][4] ), .C(\i_fifo_tx/mem[42][4] ), .D(
        \i_fifo_tx/mem[43][4] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n455 ) );
  IMUX40 \i_fifo_tx/U485  ( .A(\i_fifo_tx/mem[32][4] ), .B(
        \i_fifo_tx/mem[33][4] ), .C(\i_fifo_tx/mem[34][4] ), .D(
        \i_fifo_tx/mem[35][4] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n454 ) );
  IMUX40 \i_fifo_tx/U484  ( .A(\i_fifo_tx/mem[36][4] ), .B(
        \i_fifo_tx/mem[37][4] ), .C(\i_fifo_tx/mem[38][4] ), .D(
        \i_fifo_tx/mem[39][4] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n456 ) );
  IMUX40 \i_fifo_tx/U395  ( .A(\i_fifo_tx/n454 ), .B(\i_fifo_tx/n455 ), .C(
        \i_fifo_tx/n456 ), .D(\i_fifo_tx/n457 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n453 ) );
  IMUX40 \i_fifo_tx/U479  ( .A(\i_fifo_tx/mem[56][4] ), .B(
        \i_fifo_tx/mem[57][4] ), .C(\i_fifo_tx/mem[58][4] ), .D(
        \i_fifo_tx/mem[59][4] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n450 ) );
  IMUX40 \i_fifo_tx/U481  ( .A(\i_fifo_tx/mem[48][4] ), .B(
        \i_fifo_tx/mem[49][4] ), .C(\i_fifo_tx/mem[50][4] ), .D(
        \i_fifo_tx/mem[51][4] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n449 ) );
  IMUX40 \i_fifo_tx/U480  ( .A(\i_fifo_tx/mem[52][4] ), .B(
        \i_fifo_tx/mem[53][4] ), .C(\i_fifo_tx/mem[54][4] ), .D(
        \i_fifo_tx/mem[55][4] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n451 ) );
  IMUX40 \i_fifo_tx/U394  ( .A(\i_fifo_tx/n449 ), .B(\i_fifo_tx/n450 ), .C(
        \i_fifo_tx/n451 ), .D(\i_fifo_tx/n452 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n448 ) );
  IMUX40 \i_fifo_tx/U503  ( .A(\i_fifo_tx/mem[24][5] ), .B(
        \i_fifo_tx/mem[25][5] ), .C(\i_fifo_tx/mem[26][5] ), .D(
        \i_fifo_tx/mem[27][5] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n480 ) );
  IMUX40 \i_fifo_tx/U505  ( .A(\i_fifo_tx/mem[16][5] ), .B(
        \i_fifo_tx/mem[17][5] ), .C(\i_fifo_tx/mem[18][5] ), .D(
        \i_fifo_tx/mem[19][5] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n479 ) );
  IMUX40 \i_fifo_tx/U504  ( .A(\i_fifo_tx/mem[20][5] ), .B(
        \i_fifo_tx/mem[21][5] ), .C(\i_fifo_tx/mem[22][5] ), .D(
        \i_fifo_tx/mem[23][5] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n481 ) );
  IMUX40 \i_fifo_tx/U401  ( .A(\i_fifo_tx/n479 ), .B(\i_fifo_tx/n480 ), .C(
        \i_fifo_tx/n481 ), .D(\i_fifo_tx/n482 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n478 ) );
  IMUX40 \i_fifo_tx/U507  ( .A(\i_fifo_tx/mem[8][5] ), .B(
        \i_fifo_tx/mem[9][5] ), .C(\i_fifo_tx/mem[10][5] ), .D(
        \i_fifo_tx/mem[11][5] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n485 ) );
  IMUX40 \i_fifo_tx/U509  ( .A(\i_fifo_tx/mem[0][5] ), .B(
        \i_fifo_tx/mem[1][5] ), .C(\i_fifo_tx/mem[2][5] ), .D(
        \i_fifo_tx/mem[3][5] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n484 ) );
  IMUX40 \i_fifo_tx/U508  ( .A(\i_fifo_tx/mem[4][5] ), .B(
        \i_fifo_tx/mem[5][5] ), .C(\i_fifo_tx/mem[6][5] ), .D(
        \i_fifo_tx/mem[7][5] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n486 ) );
  IMUX40 \i_fifo_tx/U402  ( .A(\i_fifo_tx/n484 ), .B(\i_fifo_tx/n485 ), .C(
        \i_fifo_tx/n486 ), .D(\i_fifo_tx/n487 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n483 ) );
  IMUX40 \i_fifo_tx/U499  ( .A(\i_fifo_tx/mem[40][5] ), .B(
        \i_fifo_tx/mem[41][5] ), .C(\i_fifo_tx/mem[42][5] ), .D(
        \i_fifo_tx/mem[43][5] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n475 ) );
  IMUX40 \i_fifo_tx/U501  ( .A(\i_fifo_tx/mem[32][5] ), .B(
        \i_fifo_tx/mem[33][5] ), .C(\i_fifo_tx/mem[34][5] ), .D(
        \i_fifo_tx/mem[35][5] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n474 ) );
  IMUX40 \i_fifo_tx/U500  ( .A(\i_fifo_tx/mem[36][5] ), .B(
        \i_fifo_tx/mem[37][5] ), .C(\i_fifo_tx/mem[38][5] ), .D(
        \i_fifo_tx/mem[39][5] ), .S0(\i_fifo_tx/N30 ), .S1(n326), .Q(
        \i_fifo_tx/n476 ) );
  IMUX40 \i_fifo_tx/U400  ( .A(\i_fifo_tx/n474 ), .B(\i_fifo_tx/n475 ), .C(
        \i_fifo_tx/n476 ), .D(\i_fifo_tx/n477 ), .S0(n270), .S1(n1941), .Q(
        \i_fifo_tx/n473 ) );
  IMUX40 \i_fifo_tx/U495  ( .A(\i_fifo_tx/mem[56][5] ), .B(
        \i_fifo_tx/mem[57][5] ), .C(\i_fifo_tx/mem[58][5] ), .D(
        \i_fifo_tx/mem[59][5] ), .S0(\i_fifo_tx/N30 ), .S1(n327), .Q(
        \i_fifo_tx/n470 ) );
  IMUX40 \i_fifo_tx/U497  ( .A(\i_fifo_tx/mem[48][5] ), .B(
        \i_fifo_tx/mem[49][5] ), .C(\i_fifo_tx/mem[50][5] ), .D(
        \i_fifo_tx/mem[51][5] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n469 ) );
  IMUX40 \i_fifo_tx/U496  ( .A(\i_fifo_tx/mem[52][5] ), .B(
        \i_fifo_tx/mem[53][5] ), .C(\i_fifo_tx/mem[54][5] ), .D(
        \i_fifo_tx/mem[55][5] ), .S0(\i_fifo_tx/N30 ), .S1(n327), .Q(
        \i_fifo_tx/n471 ) );
  IMUX40 \i_fifo_tx/U399  ( .A(\i_fifo_tx/n469 ), .B(\i_fifo_tx/n470 ), .C(
        \i_fifo_tx/n471 ), .D(\i_fifo_tx/n472 ), .S0(\i_fifo_tx/N33 ), .S1(
        \i_fifo_tx/N32 ), .Q(\i_fifo_tx/n468 ) );
  IMUX40 \i_fifo_tx/U463  ( .A(\i_fifo_tx/mem[56][3] ), .B(
        \i_fifo_tx/mem[57][3] ), .C(\i_fifo_tx/mem[58][3] ), .D(
        \i_fifo_tx/mem[59][3] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n430 ) );
  IMUX40 \i_fifo_tx/U465  ( .A(\i_fifo_tx/mem[48][3] ), .B(
        \i_fifo_tx/mem[49][3] ), .C(\i_fifo_tx/mem[50][3] ), .D(
        \i_fifo_tx/mem[51][3] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n429 ) );
  IMUX40 \i_fifo_tx/U464  ( .A(\i_fifo_tx/mem[52][3] ), .B(
        \i_fifo_tx/mem[53][3] ), .C(\i_fifo_tx/mem[54][3] ), .D(
        \i_fifo_tx/mem[55][3] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n431 ) );
  IMUX40 \i_fifo_tx/U389  ( .A(\i_fifo_tx/n429 ), .B(\i_fifo_tx/n430 ), .C(
        \i_fifo_tx/n431 ), .D(\i_fifo_tx/n432 ), .S0(\i_fifo_tx/N33 ), .S1(
        \i_fifo_tx/N32 ), .Q(\i_fifo_tx/n428 ) );
  IMUX40 \i_fifo_tx/U472  ( .A(\i_fifo_tx/mem[20][3] ), .B(
        \i_fifo_tx/mem[21][3] ), .C(\i_fifo_tx/mem[22][3] ), .D(
        \i_fifo_tx/mem[23][3] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n441 ) );
  IMUX40 \i_fifo_tx/U473  ( .A(\i_fifo_tx/mem[16][3] ), .B(
        \i_fifo_tx/mem[17][3] ), .C(\i_fifo_tx/mem[18][3] ), .D(
        \i_fifo_tx/mem[19][3] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n439 ) );
  IMUX40 \i_fifo_tx/U471  ( .A(\i_fifo_tx/mem[24][3] ), .B(
        \i_fifo_tx/mem[25][3] ), .C(\i_fifo_tx/mem[26][3] ), .D(
        \i_fifo_tx/mem[27][3] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n440 ) );
  IMUX40 \i_fifo_tx/U470  ( .A(\i_fifo_tx/mem[28][3] ), .B(
        \i_fifo_tx/mem[29][3] ), .C(\i_fifo_tx/mem[30][3] ), .D(
        \i_fifo_tx/mem[31][3] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n442 ) );
  IMUX40 \i_fifo_tx/U476  ( .A(\i_fifo_tx/mem[4][3] ), .B(
        \i_fifo_tx/mem[5][3] ), .C(\i_fifo_tx/mem[6][3] ), .D(
        \i_fifo_tx/mem[7][3] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n446 ) );
  IMUX40 \i_fifo_tx/U477  ( .A(\i_fifo_tx/mem[0][3] ), .B(
        \i_fifo_tx/mem[1][3] ), .C(\i_fifo_tx/mem[2][3] ), .D(
        \i_fifo_tx/mem[3][3] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n444 ) );
  IMUX40 \i_fifo_tx/U475  ( .A(\i_fifo_tx/mem[8][3] ), .B(
        \i_fifo_tx/mem[9][3] ), .C(\i_fifo_tx/mem[10][3] ), .D(
        \i_fifo_tx/mem[11][3] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n445 ) );
  IMUX40 \i_fifo_tx/U474  ( .A(\i_fifo_tx/mem[12][3] ), .B(
        \i_fifo_tx/mem[13][3] ), .C(\i_fifo_tx/mem[14][3] ), .D(
        \i_fifo_tx/mem[15][3] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n447 ) );
  IMUX40 \i_fifo_tx/U468  ( .A(\i_fifo_tx/mem[36][3] ), .B(
        \i_fifo_tx/mem[37][3] ), .C(\i_fifo_tx/mem[38][3] ), .D(
        \i_fifo_tx/mem[39][3] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n436 ) );
  IMUX40 \i_fifo_tx/U469  ( .A(\i_fifo_tx/mem[32][3] ), .B(
        \i_fifo_tx/mem[33][3] ), .C(\i_fifo_tx/mem[34][3] ), .D(
        \i_fifo_tx/mem[35][3] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n434 ) );
  IMUX40 \i_fifo_tx/U467  ( .A(\i_fifo_tx/mem[40][3] ), .B(
        \i_fifo_tx/mem[41][3] ), .C(\i_fifo_tx/mem[42][3] ), .D(
        \i_fifo_tx/mem[43][3] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n435 ) );
  IMUX40 \i_fifo_tx/U466  ( .A(\i_fifo_tx/mem[44][3] ), .B(
        \i_fifo_tx/mem[45][3] ), .C(\i_fifo_tx/mem[46][3] ), .D(
        \i_fifo_tx/mem[47][3] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n437 ) );
  IMUX40 \i_fifo_tx/U454  ( .A(\i_fifo_tx/mem[28][2] ), .B(
        \i_fifo_tx/mem[29][2] ), .C(\i_fifo_tx/mem[30][2] ), .D(
        \i_fifo_tx/mem[31][2] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n422 ) );
  IMUX40 \i_fifo_tx/U458  ( .A(\i_fifo_tx/mem[12][2] ), .B(
        \i_fifo_tx/mem[13][2] ), .C(\i_fifo_tx/mem[14][2] ), .D(
        \i_fifo_tx/mem[15][2] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n427 ) );
  IMUX40 \i_fifo_tx/U450  ( .A(\i_fifo_tx/mem[44][2] ), .B(
        \i_fifo_tx/mem[45][2] ), .C(\i_fifo_tx/mem[46][2] ), .D(
        \i_fifo_tx/mem[47][2] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n417 ) );
  IMUX40 \i_fifo_tx/U446  ( .A(\i_fifo_tx/mem[60][2] ), .B(
        \i_fifo_tx/mem[61][2] ), .C(\i_fifo_tx/mem[62][2] ), .D(
        \i_fifo_tx/mem[63][2] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n412 ) );
  IMUX40 \i_fifo_tx/U422  ( .A(\i_fifo_tx/mem[28][0] ), .B(
        \i_fifo_tx/mem[29][0] ), .C(\i_fifo_tx/mem[30][0] ), .D(
        \i_fifo_tx/mem[31][0] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n382 ) );
  IMUX40 \i_fifo_tx/U426  ( .A(\i_fifo_tx/mem[12][0] ), .B(
        \i_fifo_tx/mem[13][0] ), .C(\i_fifo_tx/mem[14][0] ), .D(
        \i_fifo_tx/mem[15][0] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n387 ) );
  IMUX40 \i_fifo_tx/U418  ( .A(\i_fifo_tx/mem[44][0] ), .B(
        \i_fifo_tx/mem[45][0] ), .C(\i_fifo_tx/mem[46][0] ), .D(
        \i_fifo_tx/mem[47][0] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n377 ) );
  IMUX40 \i_fifo_tx/U414  ( .A(\i_fifo_tx/mem[60][0] ), .B(
        \i_fifo_tx/mem[61][0] ), .C(\i_fifo_tx/mem[62][0] ), .D(
        \i_fifo_tx/mem[63][0] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n372 ) );
  IMUX40 \i_fifo_tx/U438  ( .A(\i_fifo_tx/mem[28][1] ), .B(
        \i_fifo_tx/mem[29][1] ), .C(\i_fifo_tx/mem[30][1] ), .D(
        \i_fifo_tx/mem[31][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n402 ) );
  IMUX40 \i_fifo_tx/U442  ( .A(\i_fifo_tx/mem[12][1] ), .B(
        \i_fifo_tx/mem[13][1] ), .C(\i_fifo_tx/mem[14][1] ), .D(
        \i_fifo_tx/mem[15][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n407 ) );
  IMUX40 \i_fifo_tx/U434  ( .A(\i_fifo_tx/mem[44][1] ), .B(
        \i_fifo_tx/mem[45][1] ), .C(\i_fifo_tx/mem[46][1] ), .D(
        \i_fifo_tx/mem[47][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n397 ) );
  IMUX40 \i_fifo_tx/U430  ( .A(\i_fifo_tx/mem[60][1] ), .B(
        \i_fifo_tx/mem[61][1] ), .C(\i_fifo_tx/mem[62][1] ), .D(
        \i_fifo_tx/mem[63][1] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n392 ) );
  IMUX40 \i_fifo_tx/U527  ( .A(\i_fifo_tx/mem[56][7] ), .B(
        \i_fifo_tx/mem[57][7] ), .C(\i_fifo_tx/mem[58][7] ), .D(
        \i_fifo_tx/mem[59][7] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n510 ) );
  IMUX40 \i_fifo_tx/U528  ( .A(\i_fifo_tx/mem[52][7] ), .B(
        \i_fifo_tx/mem[53][7] ), .C(\i_fifo_tx/mem[54][7] ), .D(
        \i_fifo_tx/mem[55][7] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n511 ) );
  IMUX40 \i_fifo_tx/U529  ( .A(\i_fifo_tx/mem[48][7] ), .B(
        \i_fifo_tx/mem[49][7] ), .C(\i_fifo_tx/mem[50][7] ), .D(
        \i_fifo_tx/mem[51][7] ), .S0(n324), .S1(n328), .Q(\i_fifo_tx/n509 ) );
  IMUX40 \i_fifo_tx/U409  ( .A(\i_fifo_tx/n509 ), .B(\i_fifo_tx/n510 ), .C(
        \i_fifo_tx/n511 ), .D(\i_fifo_tx/n512 ), .S0(\i_fifo_tx/N33 ), .S1(
        \i_fifo_tx/N32 ), .Q(\i_fifo_tx/n508 ) );
  IMUX40 \i_fifo_tx/U536  ( .A(\i_fifo_tx/mem[20][7] ), .B(
        \i_fifo_tx/mem[21][7] ), .C(\i_fifo_tx/mem[22][7] ), .D(
        \i_fifo_tx/mem[23][7] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n521 ) );
  IMUX40 \i_fifo_tx/U537  ( .A(\i_fifo_tx/mem[16][7] ), .B(
        \i_fifo_tx/mem[17][7] ), .C(\i_fifo_tx/mem[18][7] ), .D(
        \i_fifo_tx/mem[19][7] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n519 ) );
  IMUX40 \i_fifo_tx/U535  ( .A(\i_fifo_tx/mem[24][7] ), .B(
        \i_fifo_tx/mem[25][7] ), .C(\i_fifo_tx/mem[26][7] ), .D(
        \i_fifo_tx/mem[27][7] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n520 ) );
  IMUX40 \i_fifo_tx/U534  ( .A(\i_fifo_tx/mem[28][7] ), .B(
        \i_fifo_tx/mem[29][7] ), .C(\i_fifo_tx/mem[30][7] ), .D(
        \i_fifo_tx/mem[31][7] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n522 ) );
  IMUX40 \i_fifo_tx/U540  ( .A(\i_fifo_tx/mem[4][7] ), .B(
        \i_fifo_tx/mem[5][7] ), .C(\i_fifo_tx/mem[6][7] ), .D(
        \i_fifo_tx/mem[7][7] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n526 ) );
  IMUX40 \i_fifo_tx/U539  ( .A(\i_fifo_tx/mem[8][7] ), .B(
        \i_fifo_tx/mem[9][7] ), .C(\i_fifo_tx/mem[10][7] ), .D(
        \i_fifo_tx/mem[11][7] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n525 ) );
  IMUX40 \i_fifo_tx/U541  ( .A(\i_fifo_tx/mem[0][7] ), .B(
        \i_fifo_tx/mem[1][7] ), .C(\i_fifo_tx/mem[2][7] ), .D(
        \i_fifo_tx/mem[3][7] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n524 ) );
  IMUX40 \i_fifo_tx/U538  ( .A(\i_fifo_tx/mem[12][7] ), .B(
        \i_fifo_tx/mem[13][7] ), .C(\i_fifo_tx/mem[14][7] ), .D(
        \i_fifo_tx/mem[15][7] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n527 ) );
  IMUX40 \i_fifo_tx/U532  ( .A(\i_fifo_tx/mem[36][7] ), .B(
        \i_fifo_tx/mem[37][7] ), .C(\i_fifo_tx/mem[38][7] ), .D(
        \i_fifo_tx/mem[39][7] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n516 ) );
  IMUX40 \i_fifo_tx/U533  ( .A(\i_fifo_tx/mem[32][7] ), .B(
        \i_fifo_tx/mem[33][7] ), .C(\i_fifo_tx/mem[34][7] ), .D(
        \i_fifo_tx/mem[35][7] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n514 ) );
  IMUX40 \i_fifo_tx/U531  ( .A(\i_fifo_tx/mem[40][7] ), .B(
        \i_fifo_tx/mem[41][7] ), .C(\i_fifo_tx/mem[42][7] ), .D(
        \i_fifo_tx/mem[43][7] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n515 ) );
  IMUX40 \i_fifo_tx/U530  ( .A(\i_fifo_tx/mem[44][7] ), .B(
        \i_fifo_tx/mem[45][7] ), .C(\i_fifo_tx/mem[46][7] ), .D(
        \i_fifo_tx/mem[47][7] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n517 ) );
  IMUX40 \i_fifo_tx/U518  ( .A(\i_fifo_tx/mem[28][6] ), .B(
        \i_fifo_tx/mem[29][6] ), .C(\i_fifo_tx/mem[30][6] ), .D(
        \i_fifo_tx/mem[31][6] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n502 ) );
  IMUX40 \i_fifo_tx/U522  ( .A(\i_fifo_tx/mem[12][6] ), .B(
        \i_fifo_tx/mem[13][6] ), .C(\i_fifo_tx/mem[14][6] ), .D(
        \i_fifo_tx/mem[15][6] ), .S0(n321), .S1(n327), .Q(\i_fifo_tx/n507 ) );
  IMUX40 \i_fifo_tx/U514  ( .A(\i_fifo_tx/mem[44][6] ), .B(
        \i_fifo_tx/mem[45][6] ), .C(\i_fifo_tx/mem[46][6] ), .D(
        \i_fifo_tx/mem[47][6] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n497 ) );
  IMUX40 \i_fifo_tx/U510  ( .A(\i_fifo_tx/mem[60][6] ), .B(
        \i_fifo_tx/mem[61][6] ), .C(\i_fifo_tx/mem[62][6] ), .D(
        \i_fifo_tx/mem[63][6] ), .S0(n321), .S1(n326), .Q(\i_fifo_tx/n492 ) );
  IMUX40 \i_fifo_tx/U486  ( .A(\i_fifo_tx/mem[28][4] ), .B(
        \i_fifo_tx/mem[29][4] ), .C(\i_fifo_tx/mem[30][4] ), .D(
        \i_fifo_tx/mem[31][4] ), .S0(\i_fifo_tx/N30 ), .S1(n328), .Q(
        \i_fifo_tx/n462 ) );
  IMUX40 \i_fifo_tx/U490  ( .A(\i_fifo_tx/mem[12][4] ), .B(
        \i_fifo_tx/mem[13][4] ), .C(\i_fifo_tx/mem[14][4] ), .D(
        \i_fifo_tx/mem[15][4] ), .S0(n321), .S1(n328), .Q(\i_fifo_tx/n467 ) );
  IMUX40 \i_fifo_tx/U482  ( .A(\i_fifo_tx/mem[44][4] ), .B(
        \i_fifo_tx/mem[45][4] ), .C(\i_fifo_tx/mem[46][4] ), .D(
        \i_fifo_tx/mem[47][4] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n457 ) );
  IMUX40 \i_fifo_tx/U478  ( .A(\i_fifo_tx/mem[60][4] ), .B(
        \i_fifo_tx/mem[61][4] ), .C(\i_fifo_tx/mem[62][4] ), .D(
        \i_fifo_tx/mem[63][4] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n452 ) );
  IMUX40 \i_fifo_tx/U502  ( .A(\i_fifo_tx/mem[28][5] ), .B(
        \i_fifo_tx/mem[29][5] ), .C(\i_fifo_tx/mem[30][5] ), .D(
        \i_fifo_tx/mem[31][5] ), .S0(\i_fifo_tx/N30 ), .S1(n326), .Q(
        \i_fifo_tx/n482 ) );
  IMUX40 \i_fifo_tx/U506  ( .A(\i_fifo_tx/mem[12][5] ), .B(
        \i_fifo_tx/mem[13][5] ), .C(\i_fifo_tx/mem[14][5] ), .D(
        \i_fifo_tx/mem[15][5] ), .S0(n324), .S1(n326), .Q(\i_fifo_tx/n487 ) );
  IMUX40 \i_fifo_tx/U498  ( .A(\i_fifo_tx/mem[44][5] ), .B(
        \i_fifo_tx/mem[45][5] ), .C(\i_fifo_tx/mem[46][5] ), .D(
        \i_fifo_tx/mem[47][5] ), .S0(\i_fifo_tx/N30 ), .S1(n327), .Q(
        \i_fifo_tx/n477 ) );
  IMUX40 \i_fifo_tx/U494  ( .A(\i_fifo_tx/mem[60][5] ), .B(
        \i_fifo_tx/mem[61][5] ), .C(\i_fifo_tx/mem[62][5] ), .D(
        \i_fifo_tx/mem[63][5] ), .S0(\i_fifo_tx/N30 ), .S1(n327), .Q(
        \i_fifo_tx/n472 ) );
  IMUX40 \i_fifo_tx/U462  ( .A(\i_fifo_tx/mem[60][3] ), .B(
        \i_fifo_tx/mem[61][3] ), .C(\i_fifo_tx/mem[62][3] ), .D(
        \i_fifo_tx/mem[63][3] ), .S0(n324), .S1(n327), .Q(\i_fifo_tx/n432 ) );
  IMUX40 \i_fifo_tx/U526  ( .A(\i_fifo_tx/mem[60][7] ), .B(
        \i_fifo_tx/mem[61][7] ), .C(\i_fifo_tx/mem[62][7] ), .D(
        \i_fifo_tx/mem[63][7] ), .S0(\i_fifo_tx/N30 ), .S1(n328), .Q(
        \i_fifo_tx/n512 ) );
  IMUX40 \i_fifo_rx/U396  ( .A(\i_fifo_rx/n389 ), .B(\i_fifo_rx/n390 ), .C(
        \i_fifo_rx/n391 ), .D(\i_fifo_rx/n392 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n388 ) );
  IMUX40 \i_fifo_rx/U401  ( .A(\i_fifo_rx/n409 ), .B(\i_fifo_rx/n410 ), .C(
        \i_fifo_rx/n411 ), .D(\i_fifo_rx/n412 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n408 ) );
  IMUX40 \i_fifo_rx/U406  ( .A(\i_fifo_rx/n429 ), .B(\i_fifo_rx/n430 ), .C(
        \i_fifo_rx/n431 ), .D(\i_fifo_rx/n432 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n428 ) );
  IMUX40 \i_fifo_rx/U411  ( .A(\i_fifo_rx/n449 ), .B(\i_fifo_rx/n450 ), .C(
        \i_fifo_rx/n451 ), .D(\i_fifo_rx/n452 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n448 ) );
  IMUX40 \i_fifo_rx/U416  ( .A(\i_fifo_rx/n469 ), .B(\i_fifo_rx/n470 ), .C(
        \i_fifo_rx/n471 ), .D(\i_fifo_rx/n472 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n468 ) );
  IMUX40 \i_fifo_rx/U421  ( .A(\i_fifo_rx/n489 ), .B(\i_fifo_rx/n490 ), .C(
        \i_fifo_rx/n491 ), .D(\i_fifo_rx/n492 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n488 ) );
  IMUX40 \i_fifo_rx/U426  ( .A(\i_fifo_rx/n509 ), .B(\i_fifo_rx/n510 ), .C(
        \i_fifo_rx/n511 ), .D(\i_fifo_rx/n512 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n508 ) );
  IMUX40 \i_fifo_rx/U431  ( .A(\i_fifo_rx/n529 ), .B(\i_fifo_rx/n530 ), .C(
        \i_fifo_rx/n531 ), .D(\i_fifo_rx/n532 ), .S0(n272), .S1(n1939), .Q(
        \i_fifo_rx/n528 ) );
  ADD21 \i_fifo_rx/add_139/U1_1_3  ( .A(n272), .B(\i_fifo_rx/add_139/carry [3]), .CO(\i_fifo_rx/add_139/carry [4]), .S(\i_fifo_rx/N691 ) );
  ADD21 \i_fifo_tx/add_180/U1_1_3  ( .A(n270), .B(\i_fifo_tx/add_180/carry [3]), .CO(\i_fifo_tx/add_180/carry [4]), .S(\i_fifo_tx/N158 ) );
  XOR31 \i_cordic/S1/add_53/U1_5  ( .A(\i_cordic/cor_y_s0[1][5] ), .B(
        \i_cordic/cor_x_s0[1][5] ), .C(\i_cordic/S1/add_53/carry [5]), .Q(
        \i_cordic/S1/N26 ) );
  ADD31 \i_cordic/S1/add_50/U1_4  ( .A(\i_cordic/cor_x_s0[1][4] ), .B(
        \i_cordic/cor_y_s0[1][5] ), .CI(\i_cordic/S1/add_50/carry [4]), .CO(
        \i_cordic/S1/add_50/carry [5]), .S(\i_cordic/S1/N7 ) );
  XOR31 \i_cordic/S1/add_50/U1_5  ( .A(\i_cordic/cor_x_s0[1][5] ), .B(
        \i_cordic/cor_y_s0[1][5] ), .C(\i_cordic/S1/add_50/carry [5]), .Q(
        \i_cordic/S1/N8 ) );
  ADD31 \i_cordic/S1/add_53/U1_1  ( .A(\i_cordic/cor_y_s0[1][1] ), .B(
        \i_cordic/cor_x_s0[1][2] ), .CI(\i_cordic/S1/add_53/carry [1]), .CO(
        \i_cordic/S1/add_53/carry [2]), .S(\i_cordic/S1/N22 ) );
  ADD31 \i_cordic/S1/add_50/U1_2  ( .A(\i_cordic/cor_x_s0[1][2] ), .B(
        \i_cordic/cor_y_s0[1][3] ), .CI(\i_cordic/S1/add_50/carry [2]), .CO(
        \i_cordic/S1/add_50/carry [3]), .S(\i_cordic/S1/N5 ) );
  ADD31 \i_cordic/S1/add_53/U1_2  ( .A(\i_cordic/cor_y_s0[1][2] ), .B(
        \i_cordic/cor_x_s0[1][3] ), .CI(\i_cordic/S1/add_53/carry [2]), .CO(
        \i_cordic/S1/add_53/carry [3]), .S(\i_cordic/S1/N23 ) );
  ADD31 \i_cordic/S1/add_50/U1_3  ( .A(\i_cordic/cor_x_s0[1][3] ), .B(
        \i_cordic/cor_y_s0[1][4] ), .CI(\i_cordic/S1/add_50/carry [3]), .CO(
        \i_cordic/S1/add_50/carry [4]), .S(\i_cordic/S1/N6 ) );
  DFEC3 \i_fifo_rx/wr_ptr_reg[5]  ( .D(\i_fifo_rx/N85 ), .E(\i_fifo_rx/n171 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/N38 ), .QN(\i_fifo_rx/n47 ) );
  DFEC3 \i_fifo_tx/wr_ptr_reg[5]  ( .D(\i_fifo_tx/N133 ), .E(\i_fifo_tx/n152 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/N29 ), .QN(\i_fifo_tx/n172 )
         );
  LOGIC1 U150 ( .Q(\*Logic1* ) );
  MUX22 U158 ( .A(n44), .B(n83), .S(\i_fifo_tx/n153 ), .Q(n114) );
  IMUX40 U159 ( .A(\i_fifo_tx/n243 ), .B(\i_fifo_tx/n233 ), .C(
        \i_fifo_tx/n238 ), .D(\i_fifo_tx/n228 ), .S0(\i_fifo_tx/N29 ), .S1(
        \i_fifo_tx/N28 ), .Q(n83) );
  MUX22 U160 ( .A(n45), .B(n84), .S(\i_fifo_tx/n153 ), .Q(n124) );
  IMUX40 U161 ( .A(\i_fifo_tx/n223 ), .B(\i_fifo_tx/n213 ), .C(
        \i_fifo_tx/n218 ), .D(\i_fifo_tx/n208 ), .S0(\i_fifo_tx/N29 ), .S1(
        \i_fifo_tx/N28 ), .Q(n84) );
  MUX22 U166 ( .A(\i_cordic/qbb_ibuff [2]), .B(\i_cordic/N8 ), .S(
        \i_cordic/S0/N32 ), .Q(\i_cordic/cor_y_s0[0][2] ) );
  IMAJ31 U167 ( .A(n377), .B(n236), .C(\i_cordic/cor_x_s1[2][5] ), .Q(
        \i_cordic/S2/sub_53/carry[5] ) );
  MUX22 U168 ( .A(\i_iq_demod/filtre_Q/tot [5]), .B(
        \i_iq_demod/filtre_Q/n_temp [5]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N20 ) );
  MUX22 U169 ( .A(\i_iq_demod/filtre_I/tot [5]), .B(
        \i_iq_demod/filtre_I/n_temp [5]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N20 ) );
  IMAJ31 U180 ( .A(net43019), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[2] ), .C(n503), .Q(n501) );
  MUX22 U181 ( .A(\i_cordic/qbb_ibuff [3]), .B(\i_cordic/N9 ), .S(
        \i_cordic/S0/N32 ), .Q(\i_cordic/cor_y_s0[0][3] ) );
  IMAJ31 U182 ( .A(\i_iq_demod/filtre_Q/mult2 [10]), .B(
        \i_iq_demod/filtre_Q/mult1 [10]), .C(n1178), .Q(n1176) );
  IMAJ31 U183 ( .A(\i_iq_demod/filtre_I/mult2 [10]), .B(
        \i_iq_demod/filtre_I/mult1 [10]), .C(
        \i_iq_demod/filtre_I/tot_adder/n35 ), .Q(
        \i_iq_demod/filtre_I/tot_adder/n33 ) );
  MUX22 U184 ( .A(\i_iq_demod/filtre_Q/tot [6]), .B(
        \i_iq_demod/filtre_Q/n_temp [6]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N21 ) );
  MUX22 U185 ( .A(\i_iq_demod/filtre_I/tot [6]), .B(
        \i_iq_demod/filtre_I/n_temp [6]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N21 ) );
  IMAJ31 U187 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_0_net_[5] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[4] ), .C(n594), .Q(n592)
         );
  IMAJ31 U188 ( .A(n973), .B(\i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[4] ), .C(\i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[5] ), .Q(n971) );
  IMAJ31 U192 ( .A(n1676), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[6] ), .C(n423), .Q(n422)
         );
  XNR31 U198 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][8] ), .C(n1011), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][7] ) );
  MUX22 U201 ( .A(\i_cordic/qbb_ibuff [1]), .B(\i_cordic/N7 ), .S(
        \i_cordic/S0/N32 ), .Q(\i_cordic/cor_y_s0[0][1] ) );
  XOR31 U202 ( .A(n1143), .B(n1144), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[1] ), .Q(n1150) );
  XOR31 U203 ( .A(n764), .B(n765), .C(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[1] ), .Q(n771) );
  NOR21 U204 ( .A(\i_mod_iq/fsm_mapping/n145 ), .B(\i_mod_iq/fsm_mapping/n143 ), .Q(n85) );
  MUX22 U206 ( .A(\i_iq_demod/filtre_Q/tot [7]), .B(
        \i_iq_demod/filtre_Q/n_temp [7]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N22 ) );
  MUX22 U207 ( .A(\i_iq_demod/filtre_I/tot [7]), .B(
        \i_iq_demod/filtre_I/n_temp [7]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N22 ) );
  IMAJ31 U209 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[5] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[4] ), .C(n784), .Q(n782)
         );
  MAJ31 U213 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[9] ), .C(n585), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][8] ) );
  MAJ31 U214 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[9] ), .C(n964), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][8] ) );
  IMAJ31 U215 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[2] ), .C(n625), .Q(n623)
         );
  AOI211 U223 ( .A(n86), .B(n87), .C(n88), .Q(n349) );
  INV3 U224 ( .A(n345), .Q(n88) );
  NAND31 U225 ( .A(\i_cordic/sub_173/carry [3]), .B(\i_cordic/S0/N32 ), .C(
        n177), .Q(n89) );
  INV3 U226 ( .A(n89), .Q(n275) );
  XOR31 U227 ( .A(n1197), .B(n1150), .C(n1151), .Q(
        \i_iq_demod/filtre_Q/mult2 [13]) );
  XOR31 U228 ( .A(n1186), .B(n771), .C(n772), .Q(
        \i_iq_demod/filtre_I/mult2 [13]) );
  IMAJ31 U229 ( .A(\i_iq_demod/filtre_Q/tot [10]), .B(
        \i_iq_demod/filtre_Q/temp [10]), .C(n1251), .Q(n1249) );
  IMAJ31 U230 ( .A(\i_iq_demod/filtre_I/tot [10]), .B(
        \i_iq_demod/filtre_I/temp [10]), .C(
        \i_iq_demod/filtre_I/temp_adder/n42 ), .Q(
        \i_iq_demod/filtre_I/temp_adder/n40 ) );
  IMUX21 U231 ( .A(\i_mod_iq/fsm_mapping/temp_QBB [0]), .B(
        \i_mod_iq/fsm_mapping/n154 ), .S(\i_mod_iq/fsm_mapping/n92 ), .Q(
        \i_mod_iq/fsm_mapping/n159 ) );
  MUX22 U232 ( .A(\i_iq_demod/filtre_Q/tot [8]), .B(
        \i_iq_demod/filtre_Q/n_temp [8]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N23 ) );
  MUX22 U233 ( .A(\i_iq_demod/filtre_I/tot [8]), .B(
        \i_iq_demod/filtre_I/n_temp [8]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N23 ) );
  MAJ31 U236 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[9] ), .C(n775), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][8] ) );
  IMAJ31 U238 ( .A(n1726), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[2] ), .C(n647), .Q(n645)
         );
  MAJ31 U239 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_6_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][8] ), .C(n608), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][8] ) );
  IMAJ31 U241 ( .A(n1759), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[2] ), .C(n814), .Q(n812)
         );
  MAJ31 U243 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][8] ), .C(n987), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][8] ) );
  XNR31 U246 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][8] ), .C(n843), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][7] ) );
  XNR31 U248 ( .A(n935), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[9][4] ), .C(n1188), 
        .Q(\i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][3] ) );
  XNR31 U251 ( .A(n556), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[9][4] ), .C(
        \i_iq_demod/filtre_I/mult1_multiplier/n17 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][3] ) );
  NAND31 U252 ( .A(n99), .B(\i_cordic/cor_x_s1[2][2] ), .C(n225), .Q(n371) );
  AOI211 U253 ( .A(\i_fifo_rx/n153 ), .B(\i_fifo_rx/N40 ), .C(n346), .Q(n348)
         );
  NOR40 U254 ( .A(\i_cordic/qbb_ibuff [3]), .B(\i_cordic/qbb_ibuff [2]), .C(
        \i_cordic/qbb_ibuff [1]), .D(\i_cordic/N6 ), .Q(
        \i_cordic/sub_170/carry [4]) );
  OAI212 U257 ( .A(\i_fifo_tx/n180 ), .B(\i_fifo_tx/N31 ), .C(n336), .Q(n90)
         );
  INV3 U258 ( .A(n90), .Q(n340) );
  XNR31 U259 ( .A(\i_iq_demod/filtre_Q/mult2 [13]), .B(
        \i_iq_demod/filtre_Q/mult1 [13]), .C(n1170), .Q(
        \i_iq_demod/filtre_Q/tot [13]) );
  XNR31 U260 ( .A(\i_iq_demod/filtre_I/mult2 [13]), .B(
        \i_iq_demod/filtre_I/mult1 [13]), .C(
        \i_iq_demod/filtre_I/tot_adder/n27 ), .Q(\i_iq_demod/filtre_I/tot [13]) );
  IMUX21 U261 ( .A(\i_mod_iq/fsm_mapping/n129 ), .B(
        \i_mod_iq/fsm_mapping/S_AQ ), .S(\i_mod_iq/fsm_mapping/n92 ), .Q(
        \i_mod_iq/fsm_mapping/n132 ) );
  OAI212 U262 ( .A(\i_mod_iq/fsm_mapping/n98 ), .B(\i_mod_iq/fsm_mapping/n163 ), .C(\i_mod_iq/fsm_mapping/n69 ), .Q(\i_mod_iq/fsm_mapping/n81 ) );
  MUX22 U265 ( .A(\i_iq_demod/filtre_Q/tot [9]), .B(
        \i_iq_demod/filtre_Q/n_temp [9]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N24 ) );
  MUX22 U268 ( .A(\i_iq_demod/filtre_I/tot [9]), .B(
        \i_iq_demod/filtre_I/n_temp [9]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N24 ) );
  MAJ31 U275 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][8] ), .C(n798), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][8] ) );
  IMAJ31 U277 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_0_net_[3] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[2] ), .C(n411), .Q(n409)
         );
  MAJ31 U278 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_6_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[2][8] ), .C(n419), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][8] ) );
  XNR31 U281 ( .A(n1125), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[9][4] ), .C(n1194), 
        .Q(\i_iq_demod/filtre_Q/mult2_multiplier/register_pipe[10][3] ) );
  XNR31 U282 ( .A(n746), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register_pipe[9][4] ), .C(n1183), 
        .Q(\i_iq_demod/filtre_I/mult2_multiplier/register_pipe[10][3] ) );
  XNR31 U284 ( .A(n1056), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][8] ), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[9] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[6][7] ) );
  MUX22 U285 ( .A(\i_cordic/qbb_ibuff [4]), .B(\i_cordic/N10 ), .S(
        \i_cordic/S0/N32 ), .Q(\i_cordic/cor_y_s0[0][4] ) );
  IMAJ31 U286 ( .A(n229), .B(\i_cordic/cor_x_s1[2][4] ), .C(n373), .Q(n376) );
  IMAJ31 U288 ( .A(\i_iq_demod/filtre_Q/mult2 [2]), .B(
        \i_iq_demod/filtre_Q/mult1 [2]), .C(n1166), .Q(n1164) );
  IMAJ31 U289 ( .A(\i_iq_demod/filtre_Q/mult2 [6]), .B(
        \i_iq_demod/filtre_Q/mult1 [6]), .C(n1158), .Q(n1156) );
  XNR31 U290 ( .A(n953), .B(n954), .C(n1191), .Q(n960) );
  XNR31 U291 ( .A(n510), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[6][7] ), .C(
        \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[7] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[7][6] ) );
  IMAJ31 U292 ( .A(\i_iq_demod/filtre_I/mult2 [2]), .B(
        \i_iq_demod/filtre_I/mult1 [2]), .C(
        \i_iq_demod/filtre_I/tot_adder/n15 ), .Q(
        \i_iq_demod/filtre_I/tot_adder/n13 ) );
  IMAJ31 U293 ( .A(\i_iq_demod/filtre_I/mult2 [6]), .B(
        \i_iq_demod/filtre_I/mult1 [6]), .C(\i_iq_demod/filtre_I/tot_adder/n7 ), .Q(\i_iq_demod/filtre_I/tot_adder/n5 ) );
  XNR31 U294 ( .A(n574), .B(n575), .C(
        \i_iq_demod/filtre_I/mult1_multiplier/n20 ), .Q(n581) );
  AOI211 U295 ( .A(\i_fifo_tx/n180 ), .B(\i_fifo_tx/N31 ), .C(n337), .Q(n339)
         );
  NAND22 U296 ( .A(\i_iq_demod/sine_IN [0]), .B(\i_iq_demod/gen_sin/n2 ), .Q(
        \i_iq_demod/demod/n22 ) );
  AOI211 U297 ( .A(\i_iq_demod/demod/n32 ), .B(\i_iq_demod/demod/n33 ), .C(
        \i_iq_demod/demod/n43 ), .Q(\i_iq_demod/demod/IC [0]) );
  MUX31 U298 ( .A(\i_mod_iq/fsm_mapping/n139 ), .B(\i_mod_iq/fsm_mapping/n134 ), .C(\i_mod_iq/fsm_mapping/n134 ), .S0(\i_mod_iq/fsm_mapping/n145 ), .S1(
        \i_mod_iq/fsm_mapping/n143 ), .Q(\i_mod_iq/fsm_mapping/n140 ) );
  NAND41 U299 ( .A(fifo_rx_psel_i), .B(n37), .C(mux_i[1]), .D(\i_fifo_rx/n11 ), 
        .Q(\i_fifo_rx/n172 ) );
  MUX22 U302 ( .A(\i_iq_demod/filtre_Q/tot [11]), .B(
        \i_iq_demod/filtre_Q/n_temp [11]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N26 ) );
  MUX22 U305 ( .A(\i_iq_demod/filtre_I/tot [11]), .B(
        \i_iq_demod/filtre_I/n_temp [11]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N26 ) );
  MAJ31 U309 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_9_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][8] ), .C(n1628), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][8] ) );
  MAJ31 U311 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][8] ), .C(n821), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][8] ) );
  MAJ31 U313 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][8] ), .C(n1011), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][8] ) );
  MAJ31 U315 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_9_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][8] ), .C(n442), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][8] ) );
  IMAJ31 U316 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[6][2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[2] ), .C(n522), .Q(n520) );
  NOR21 U321 ( .A(n95), .B(n96), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_51_net_[1] ) );
  NOR31 U322 ( .A(\i_cdr/i_bit_recovery/phase_q [1]), .B(n260), .C(
        \i_cdr/i_bit_recovery/phase_q [0]), .Q(n381) );
  NOR21 U323 ( .A(n97), .B(n98), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_51_net_[1] ) );
  AOI2111 U324 ( .A(n99), .B(n218), .C(n225), .D(n100), .Q(n361) );
  XOR31 U327 ( .A(n1208), .B(\i_iq_demod/filtre_Q/data_2_1 [4]), .C(
        \i_iq_demod/filtre_Q/data_1_1 [4]), .Q(n173) );
  XOR31 U329 ( .A(n1217), .B(\i_iq_demod/filtre_Q/data_2_2 [4]), .C(
        \i_iq_demod/filtre_Q/data_1_2 [4]), .Q(n210) );
  IMAJ31 U331 ( .A(\i_iq_demod/filtre_Q/mult2 [4]), .B(
        \i_iq_demod/filtre_Q/mult1 [4]), .C(n1162), .Q(n1160) );
  IMAJ31 U332 ( .A(\i_iq_demod/filtre_Q/mult2 [8]), .B(
        \i_iq_demod/filtre_Q/mult1 [8]), .C(n1154), .Q(n1152) );
  XOR31 U333 ( .A(n1192), .B(n960), .C(n961), .Q(
        \i_iq_demod/filtre_Q/mult1 [13]) );
  IMAJ31 U336 ( .A(\i_iq_demod/filtre_I/mult2 [4]), .B(
        \i_iq_demod/filtre_I/mult1 [4]), .C(
        \i_iq_demod/filtre_I/tot_adder/n11 ), .Q(
        \i_iq_demod/filtre_I/tot_adder/n9 ) );
  IMAJ31 U337 ( .A(\i_iq_demod/filtre_I/mult2 [8]), .B(
        \i_iq_demod/filtre_I/mult1 [8]), .C(\i_iq_demod/filtre_I/tot_adder/n3 ), .Q(\i_iq_demod/filtre_I/tot_adder/n1 ) );
  XOR31 U338 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/n21 ), .B(n581), .C(
        n582), .Q(\i_iq_demod/filtre_I/mult1 [13]) );
  MUX22 U339 ( .A(\i_cordic/N6 ), .B(\i_cordic/N6 ), .S(\i_cordic/S0/N32 ), 
        .Q(\i_cordic/cor_y_s0[0][0] ) );
  NAND22 U340 ( .A(n101), .B(n329), .Q(\i_cordic/S2/sub_56/carry[5] ) );
  NOR31 U341 ( .A(demod_iq_qif_i[3]), .B(demod_iq_qif_i[2]), .C(n335), .Q(
        \i_iq_demod/demod/r70/carry [4]) );
  INV3 U343 ( .A(n102), .Q(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/carry [3]) );
  INV3 U345 ( .A(n103), .Q(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/carry [3]) );
  AOI211 U346 ( .A(\i_iq_demod/demod/n20 ), .B(\i_iq_demod/demod/n22 ), .C(
        \i_iq_demod/demod/n31 ), .Q(\i_iq_demod/demod/QS [0]) );
  MUX22 U347 ( .A(\i_mod_iq/fsm_mapping/n84 ), .B(\i_mod_iq/fsm_mapping/n89 ), 
        .S(\i_mod_iq/fsm_mapping/n92 ), .Q(\i_mod_iq/fsm_mapping/n88 ) );
  IMUX21 U349 ( .A(\i_fifo_rx/shift_register [2]), .B(\i_fifo_rx/N92 ), .S(
        \i_fifo_rx/n170 ), .Q(n106) );
  MUX22 U353 ( .A(\i_iq_demod/filtre_Q/tot [12]), .B(
        \i_iq_demod/filtre_Q/n_temp [12]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N27 ) );
  MUX22 U356 ( .A(\i_iq_demod/filtre_I/tot [12]), .B(
        \i_iq_demod/filtre_I/n_temp [12]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N27 ) );
  IMUX21 U357 ( .A(\i_mod_iq/fsm_mapping/n187 ), .B(\i_mod_iq/fsm_mapping/n65 ), .S(\i_mod_iq/fsm_mapping/n82 ), .Q(\i_mod_iq/fsm_mapping/n185 ) );
  MUX22 U359 ( .A(\i_cordic/S3/N37 ), .B(\i_cordic/S3/N37 ), .S(
        \i_cordic/S2/n21 ), .Q(\i_cordic/cor_w_s1[4][4] ) );
  XOR31 U362 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_9_net_[6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][6] ), .C(n636), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][5] ) );
  XOR31 U363 ( .A(n1015), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][6] ), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[6] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][5] ) );
  NOR31 U366 ( .A(\i_cordic/qbb_ibuff [2]), .B(\i_cordic/qbb_ibuff [1]), .C(
        \i_cordic/N6 ), .Q(\i_cordic/sub_170/carry [3]) );
  MAJ31 U368 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][8] ), .C(n843), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][8] ) );
  MAJ31 U370 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_12_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][8] ), .C(n464), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[5][8] ) );
  XOR31 U371 ( .A(n1134), .B(n1135), .C(n1196), .Q(n1144) );
  XOR31 U372 ( .A(n944), .B(n945), .C(n1190), .Q(n954) );
  XOR31 U373 ( .A(n755), .B(n756), .C(n1185), .Q(n765) );
  XOR31 U374 ( .A(n565), .B(n566), .C(
        \i_iq_demod/filtre_I/mult1_multiplier/n19 ), .Q(n575) );
  IMAJ31 U376 ( .A(\i_iq_demod/filtre_Q/data_2_1 [2]), .B(
        \i_iq_demod/filtre_Q/data_1_1 [2]), .C(n1212), .Q(n1211) );
  IMAJ31 U377 ( .A(\i_iq_demod/filtre_Q/data_2_2 [2]), .B(
        \i_iq_demod/filtre_Q/data_1_2 [2]), .C(n1767), .Q(n1220) );
  IMAJ31 U379 ( .A(n383), .B(\i_cdr/i_bit_recovery/phase_q [2]), .C(n264), .Q(
        n386) );
  OAI212 U380 ( .A(\i_cordic/S0/N32 ), .B(\i_cordic/n5 ), .C(\i_cordic/N13 ), 
        .Q(\i_cordic/n22 ) );
  NOR31 U381 ( .A(demod_iq_iif_i[3]), .B(demod_iq_iif_i[2]), .C(n334), .Q(
        \i_iq_demod/demod/r69/carry [4]) );
  IMAJ31 U383 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[8][2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[2] ), .C(n740), .Q(n738) );
  IMAJ31 U387 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[8][2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[2] ), .C(n1119), .Q(
        n1117) );
  NAND22 U388 ( .A(\i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [1]), .B(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/carry [1]), .Q(n110) );
  IMAJ31 U390 ( .A(\i_iq_demod/filtre_Q/tot [2]), .B(
        \i_iq_demod/filtre_Q/temp [2]), .C(n1240), .Q(n1238) );
  IMAJ31 U391 ( .A(\i_iq_demod/filtre_Q/tot [6]), .B(
        \i_iq_demod/filtre_Q/temp [6]), .C(n1232), .Q(n1230) );
  IMAJ31 U393 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[8][2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[2] ), .C(n550), .Q(n548) );
  NAND22 U394 ( .A(\i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [1]), .B(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/carry [1]), .Q(n111) );
  XOR31 U396 ( .A(\i_cdr/i_cdr/n8 ), .B(\i_cdr/i_cdr/n7 ), .C(
        \i_cdr/i_cdr/count [0]), .Q(n394) );
  IMAJ31 U397 ( .A(\i_iq_demod/filtre_I/tot [2]), .B(
        \i_iq_demod/filtre_I/temp [2]), .C(
        \i_iq_demod/filtre_I/temp_adder/n15 ), .Q(
        \i_iq_demod/filtre_I/temp_adder/n13 ) );
  IMAJ31 U398 ( .A(\i_iq_demod/filtre_I/tot [6]), .B(
        \i_iq_demod/filtre_I/temp [6]), .C(\i_iq_demod/filtre_I/temp_adder/n7 ), .Q(\i_iq_demod/filtre_I/temp_adder/n5 ) );
  IMUX21 U399 ( .A(\i_fifo_rx/shift_register [0]), .B(\i_fifo_rx/N94 ), .S(
        \i_fifo_rx/n170 ), .Q(n112) );
  NAND22 U401 ( .A(\i_iq_demod/demod/QS [0]), .B(\i_iq_demod/demod/IC [0]), 
        .Q(n113) );
  INV3 U402 ( .A(n113), .Q(\i_iq_demod/demod/dp_cluster_1/add_87/carry [1]) );
  MUX22 U404 ( .A(\i_iq_demod/filtre_Q/tot [10]), .B(
        \i_iq_demod/filtre_Q/n_temp [10]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N25 ) );
  IMAJ31 U405 ( .A(\i_iq_demod/filtre_Q/tot [12]), .B(
        \i_iq_demod/filtre_Q/temp [12]), .C(n1246), .Q(n1245) );
  MUX22 U407 ( .A(\i_iq_demod/filtre_I/tot [10]), .B(
        \i_iq_demod/filtre_I/n_temp [10]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N25 ) );
  IMAJ31 U408 ( .A(\i_iq_demod/filtre_I/tot [12]), .B(
        \i_iq_demod/filtre_I/temp [12]), .C(
        \i_iq_demod/filtre_I/temp_adder/n35 ), .Q(
        \i_iq_demod/filtre_I/temp_adder/n33 ) );
  IMUX21 U409 ( .A(\i_mod_iq/fsm_mapping/n147 ), .B(
        \i_mod_iq/fsm_mapping/n151 ), .S(\i_mod_iq/fsm_mapping/n92 ), .Q(
        \i_mod_iq/fsm_mapping/n148 ) );
  AOI211 U413 ( .A(\i_fifo_tx/n186 ), .B(\i_fifo_tx/N40 ), .C(n115), .Q(
        \i_fifo_tx/next_state_rd ) );
  MAJ31 U419 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][8] ), .C(n1033), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][8] ) );
  NOR31 U420 ( .A(\i_cordic/ibb_ibuff [2]), .B(\i_cordic/ibb_ibuff [1]), .C(
        \i_cordic/N13 ), .Q(\i_cordic/sub_173/carry [3]) );
  IMAJ31 U426 ( .A(n537), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[2] ), .C(
        \i_iq_demod/filtre_I/mult1_multiplier/register[7][2] ), .Q(n535) );
  NOR21 U427 ( .A(\i_cdr/i_cdr/count [3]), .B(n116), .Q(n390) );
  NAND22 U428 ( .A(\i_cordic/cor_y_s0[0][0] ), .B(\i_cordic/n22 ), .Q(
        \i_cordic/S0/sub_50/carry [1]) );
  IMAJ31 U430 ( .A(\i_iq_demod/filtre_Q/tot [4]), .B(
        \i_iq_demod/filtre_Q/temp [4]), .C(n1236), .Q(n1234) );
  IMAJ31 U431 ( .A(\i_iq_demod/filtre_Q/tot [8]), .B(
        \i_iq_demod/filtre_Q/temp [8]), .C(n1228), .Q(n1226) );
  OAI2111 U432 ( .A(n49), .B(n5), .C(\i_iq_demod/demod/validation/n5 ), .D(
        mux_i[21]), .Q(\i_iq_demod/demod/validation/n1 ) );
  XOR31 U433 ( .A(\i_cdr/i_bit_recovery/phase_q [5]), .B(n259), .C(
        \i_cdr/i_bit_recovery/sub_68/carry[5] ), .Q(
        \i_cdr/i_bit_recovery/phase_diff[5] ) );
  IMAJ31 U434 ( .A(\i_iq_demod/filtre_I/tot [4]), .B(
        \i_iq_demod/filtre_I/temp [4]), .C(
        \i_iq_demod/filtre_I/temp_adder/n11 ), .Q(
        \i_iq_demod/filtre_I/temp_adder/n9 ) );
  IMAJ31 U435 ( .A(\i_iq_demod/filtre_I/tot [8]), .B(
        \i_iq_demod/filtre_I/temp [8]), .C(\i_iq_demod/filtre_I/temp_adder/n3 ), .Q(\i_iq_demod/filtre_I/temp_adder/n1 ) );
  IMUX21 U436 ( .A(\i_fifo_rx/shift_register [1]), .B(\i_fifo_rx/N93 ), .S(
        \i_fifo_rx/n170 ), .Q(n118) );
  MAJ31 U440 ( .A(\i_iq_demod/filtre_I/data_2_2 [4]), .B(
        \i_iq_demod/filtre_I/data_1_2 [4]), .C(n1199), .Q(
        \i_iq_demod/filtre_I/_16_net_[8] ) );
  MAJ31 U442 ( .A(\i_iq_demod/filtre_Q/data_2_1 [4]), .B(
        \i_iq_demod/filtre_Q/data_1_1 [4]), .C(n1208), .Q(
        \i_iq_demod/filtre_Q/_15_net_[8] ) );
  MAJ31 U444 ( .A(\i_iq_demod/filtre_Q/data_2_2 [4]), .B(
        \i_iq_demod/filtre_Q/data_1_2 [4]), .C(n1217), .Q(
        \i_iq_demod/filtre_Q/_16_net_[8] ) );
  NAND22 U445 ( .A(\i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [3]), .B(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/carry [3]), .Q(n119) );
  XNR31 U448 ( .A(n1245), .B(\i_iq_demod/filtre_Q/tot [13]), .C(
        \i_iq_demod/filtre_Q/temp [13]), .Q(\i_iq_demod/filtre_Q/n_temp [13])
         );
  MAJ31 U450 ( .A(\i_iq_demod/filtre_I/data_2_1 [4]), .B(
        \i_iq_demod/filtre_I/data_1_1 [4]), .C(
        \i_iq_demod/filtre_I/sum1_adder/n4 ), .Q(
        \i_iq_demod/filtre_I/_15_net_[8] ) );
  NAND22 U451 ( .A(\i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [3]), .B(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/carry [3]), .Q(n120) );
  NOR21 U453 ( .A(\i_cdr/i_cdr/data_en_w ), .B(n121), .Q(\i_cdr/i_cdr/N160 )
         );
  XNR31 U455 ( .A(\i_iq_demod/filtre_I/temp_adder/n33 ), .B(
        \i_iq_demod/filtre_I/tot [13]), .C(\i_iq_demod/filtre_I/temp [13]), 
        .Q(\i_iq_demod/filtre_I/n_temp [13]) );
  NOR21 U456 ( .A(n122), .B(n123), .Q(\i_mod_iq/en_gen_map/n1 ) );
  NOR40 U458 ( .A(\i_fifo_rx/i [0]), .B(\i_fifo_rx/i [1]), .C(\i_fifo_rx/n188 ), .D(\i_fifo_rx/i [2]), .Q(\i_fifo_rx/n177 ) );
  AOI311 U462 ( .A(fifo_tx_enable_o), .B(\i_fifo_tx/state_rd ), .C(
        \i_fifo_tx/n191 ), .D(\i_fifo_tx/n78 ), .Q(n125) );
  INV3 U463 ( .A(n125), .Q(\i_fifo_tx/n204 ) );
  INV3 U464 ( .A(\i_iq_demod/filtre_I/factor/n4 ), .Q(
        \i_iq_demod/filtre_I/factor/n23 ) );
  INV3 U465 ( .A(n1263), .Q(n1274) );
  INV3 U466 ( .A(\i_iq_demod/filtre_I/_16_net_[8] ), .Q(n1187) );
  INV3 U467 ( .A(\i_iq_demod/filtre_Q/_15_net_[8] ), .Q(n1193) );
  INV3 U468 ( .A(\i_iq_demod/filtre_Q/_16_net_[8] ), .Q(n1198) );
  NAND22 U474 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/A_pipe [0]), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/B_pipe ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/n21 ) );
  NAND22 U475 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/A_pipe [0]), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/B_pipe ), .Q(n1186) );
  NAND22 U476 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/A_pipe [0]), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/B_pipe ), .Q(n1192) );
  NAND22 U477 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/A_pipe [0]), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/B_pipe ), .Q(n1197) );
  INV3 U478 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_15_net_[0] ), .Q(n507)
         );
  INV3 U480 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[0] ), .Q(n886)
         );
  XOR21 U486 ( .A(n1211), .B(n1210), .Q(n167) );
  INV3 U488 ( .A(\i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/S1/sub_50/B_not [5])
         );
  XOR21 U493 ( .A(n1202), .B(n1201), .Q(n205) );
  XNR21 U495 ( .A(\i_fifo_rx/add_90/carry [7]), .B(\i_fifo_rx/i [7]), .Q(n238)
         );
  XNR21 U496 ( .A(\i_fifo_tx/r80/carry [4]), .B(\i_fifo_tx/counter_clock [4]), 
        .Q(n245) );
  XNR21 U497 ( .A(\i_cdr/i_cdr/add_119/carry [4]), .B(\i_cdr/i_cdr/count [4]), 
        .Q(n246) );
  CLKIN0 U508 ( .A(\i_iq_demod/filtre_Q/shift_r/N3 ), .Q(n265) );
  CLKIN0 U510 ( .A(\i_iq_demod/filtre_I/shift_r/N3 ), .Q(n267) );
  NAND22 U516 ( .A(N12), .B(n71), .Q(n14) );
  INV3 U518 ( .A(\i_cdr/i_bit_recovery/n10 ), .Q(\i_cdr/i_bit_recovery/N91 )
         );
  INV3 U522 ( .A(n71), .Q(n5) );
  CLKIN1 U523 ( .A(\i_iq_demod/filtre_I/n22 ), .Q(\i_iq_demod/filtre_I/N123 )
         );
  NAND22 U524 ( .A(\i_iq_demod/filtre_I/n42 ), .B(
        \i_iq_demod/filtre_I/shift_count [1]), .Q(\i_iq_demod/filtre_I/n22 )
         );
  CLKIN1 U525 ( .A(n1391), .Q(\i_iq_demod/filtre_Q/N123 ) );
  NAND22 U526 ( .A(n1398), .B(\i_iq_demod/filtre_Q/shift_count [1]), .Q(n1391)
         );
  INV3 U535 ( .A(n289), .Q(\i_iq_demod/filtre_Q/out_factor1_req [1]) );
  INV3 U536 ( .A(n290), .Q(\i_iq_demod/filtre_I/out_factor1_req [1]) );
  INV3 U537 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_0_net_[6] ), .Q(n583)
         );
  INV3 U538 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[6] ), .Q(n773)
         );
  INV3 U539 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[6] ), .Q(n962)
         );
  INV3 U540 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_0_net_[6] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/genblk1[0].adder/n10 ) );
  NOR21 U542 ( .A(\i_cordic/ibb_ibuff [1]), .B(\i_cordic/N13 ), .Q(
        \i_cordic/sub_173/carry [2]) );
  NOR21 U543 ( .A(\i_cordic/qbb_ibuff [1]), .B(\i_cordic/N6 ), .Q(
        \i_cordic/sub_170/carry [2]) );
  XOR21 U551 ( .A(\i_cordic/sub_173/carry [2]), .B(n178), .Q(\i_cordic/N15 )
         );
  XOR21 U552 ( .A(\i_cordic/sub_170/carry [2]), .B(\i_cordic/n12 ), .Q(
        \i_cordic/N8 ) );
  XOR21 U553 ( .A(\i_cordic/sub_173/carry [3]), .B(n177), .Q(\i_cordic/N16 )
         );
  XOR21 U554 ( .A(\i_cordic/sub_170/carry [3]), .B(\i_cordic/n10 ), .Q(
        \i_cordic/N9 ) );
  INV3 U555 ( .A(n331), .Q(\i_cordic/S0/sub_53/carry [1]) );
  NOR21 U556 ( .A(\i_cordic/n22 ), .B(\i_cordic/cor_y_s0[0][0] ), .Q(n331) );
  XOR21 U557 ( .A(n179), .B(n213), .Q(\i_cordic/N14 ) );
  XOR21 U558 ( .A(\i_cordic/n16 ), .B(\i_cordic/n14 ), .Q(\i_cordic/N7 ) );
  NOR21 U559 ( .A(\i_cordic/S0/sub_50/B_not [0]), .B(\i_cordic/n22 ), .Q(
        \i_cordic/S0/r64/carry [1]) );
  XNR21 U560 ( .A(\i_cordic/qbb_ibuff [4]), .B(\i_cordic/sub_170/carry [4]), 
        .Q(\i_cordic/N10 ) );
  NOR21 U561 ( .A(demod_iq_qif_i[2]), .B(n335), .Q(
        \i_iq_demod/demod/r70/carry [3]) );
  INV3 U562 ( .A(\i_iq_demod/demod/r70/carry [2]), .Q(n335) );
  NOR21 U563 ( .A(demod_iq_qif_i[1]), .B(\i_iq_demod/demod/N41 ), .Q(
        \i_iq_demod/demod/r70/carry [2]) );
  NOR21 U564 ( .A(\i_iq_demod/gen_sin/next_state [0]), .B(
        \i_iq_demod/gen_sin/current_state [2]), .Q(\i_iq_demod/gen_sin/n6 ) );
  NOR21 U565 ( .A(demod_iq_iif_i[1]), .B(\i_iq_demod/demod/N36 ), .Q(
        \i_iq_demod/demod/r69/carry [2]) );
  NOR21 U566 ( .A(demod_iq_iif_i[2]), .B(n334), .Q(
        \i_iq_demod/demod/r69/carry [3]) );
  INV3 U567 ( .A(\i_iq_demod/demod/r69/carry [2]), .Q(n334) );
  NOR21 U568 ( .A(n1384), .B(n1385), .Q(\i_iq_demod/filtre_Q/sel [2]) );
  NOR21 U569 ( .A(\i_cdr/i_cdr/n7 ), .B(\i_cdr/i_cdr/curr_state[1] ), .Q(
        \i_cdr/i_cdr/cycles[2] ) );
  NOR31 U570 ( .A(\i_iq_demod/gen_sin/current_state [2]), .B(
        \i_iq_demod/gen_sin/n2 ), .C(\i_iq_demod/gen_sin/current_state [0]), 
        .Q(\i_iq_demod/cosine_IN [1]) );
  NOR21 U571 ( .A(\i_iq_demod/filtre_I/n1 ), .B(\i_iq_demod/filtre_I/n2 ), .Q(
        \i_iq_demod/filtre_I/sel [2]) );
  NOR21 U572 ( .A(\i_mod_iq/fsm_mapping/n214 ), .B(\i_mod_iq/fsm_mapping/n215 ), .Q(\i_mod_iq/fsm_mapping/n173 ) );
  XNR21 U587 ( .A(\i_cordic/cor_x_s0[0][0] ), .B(\i_cordic/S0/sub_50/B_not [0]), .Q(\i_cordic/S0/N9 ) );
  XNR21 U588 ( .A(\i_cordic/cor_x_s0[0][0] ), .B(\i_cordic/cor_y_s0[0][0] ), 
        .Q(n276) );
  NOR21 U591 ( .A(\i_cordic/S2/N29 ), .B(\i_cordic/S2/N30 ), .Q(n329) );
  INV3 U598 ( .A(N12), .Q(N13) );
  INV3 U599 ( .A(N10), .Q(N11) );
  XOR21 U600 ( .A(demod_iq_qif_i[4]), .B(\i_iq_demod/demod/r70/carry [4]), .Q(
        n278) );
  XNR21 U601 ( .A(\i_iq_demod/demod/r70/carry [3]), .B(\i_iq_demod/demod/n25 ), 
        .Q(n279) );
  XNR21 U602 ( .A(\i_iq_demod/demod/r70/carry [2]), .B(\i_iq_demod/demod/n27 ), 
        .Q(n280) );
  XNR21 U603 ( .A(\i_iq_demod/demod/n31 ), .B(\i_iq_demod/demod/n29 ), .Q(n281) );
  XNR21 U604 ( .A(\i_iq_demod/demod/n43 ), .B(\i_iq_demod/demod/n41 ), .Q(n282) );
  XNR21 U605 ( .A(\i_iq_demod/demod/r69/carry [2]), .B(\i_iq_demod/demod/n39 ), 
        .Q(n283) );
  XNR21 U606 ( .A(\i_iq_demod/demod/r69/carry [3]), .B(\i_iq_demod/demod/n37 ), 
        .Q(n284) );
  XOR21 U607 ( .A(demod_iq_iif_i[4]), .B(\i_iq_demod/demod/r69/carry [4]), .Q(
        n285) );
  NAND22 U608 ( .A(\i_iq_demod/demod/validation/n2 ), .B(
        \i_iq_demod/demod/validation/current_state_valid [0]), .Q(
        \i_iq_demod/demod/validation/n3 ) );
  NAND22 U609 ( .A(\i_cdr/i_bit_recovery/n14 ), .B(cdr_valid_i), .Q(
        \i_cdr/i_bit_recovery/n11 ) );
  NAND22 U610 ( .A(\i_cdr/i_bit_recovery/n12 ), .B(
        \i_cdr/i_bit_recovery/curr_state [0]), .Q(\i_cdr/i_bit_recovery/n10 )
         );
  NAND22 U611 ( .A(\i_iq_demod/gen_sin/n5 ), .B(
        \i_iq_demod/gen_sin/current_state [0]), .Q(\i_iq_demod/gen_sin/n1 ) );
  NAND22 U612 ( .A(\i_fifo_tx/N144 ), .B(\i_fifo_tx/state_rd ), .Q(n286) );
  INV3 U613 ( .A(\i_mod_iq/fsm_mapping/n199 ), .Q(\i_mod_iq/fsm_mapping/n165 )
         );
  XOR21 U615 ( .A(\i_cordic/S0/n39 ), .B(\i_cordic/S0/sub_50/carry [5]), .Q(
        \i_cordic/S0/N14 ) );
  INV3 U616 ( .A(n330), .Q(\i_cordic/S1/sub_53/carry [1]) );
  NOR21 U618 ( .A(n360), .B(n333), .Q(\i_cordic/S1/add_53/carry [1]) );
  INV3 U619 ( .A(\i_cordic/cor_y_s0[1][0] ), .Q(n333) );
  XOR21 U620 ( .A(\i_cordic/cor_y_s0[0][0] ), .B(\i_cordic/n22 ), .Q(n287) );
  XNR21 U622 ( .A(\i_cordic/S2/N30 ), .B(\i_cordic/S2/N29 ), .Q(
        \i_cordic/S2/N36 ) );
  XNR21 U624 ( .A(\i_cordic/S2/sub_56/carry[5] ), .B(\i_cordic/S2/N32 ), .Q(
        \i_cordic/S2/N38 ) );
  INV3 U626 ( .A(n332), .Q(\i_iq_demod/demod/dp_cluster_0/sub_88/carry [1]) );
  NOR21 U627 ( .A(\i_iq_demod/demod/dp_cluster_0/sub_88/B_not [0]), .B(
        \i_iq_demod/demod/QC [0]), .Q(n332) );
  XOR21 U631 ( .A(\i_iq_demod/demod/dp_cluster_0/sub_mult_88/carry [1]), .B(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [1]), .Q(
        \i_iq_demod/Q_BB_IN [1]) );
  XNR21 U632 ( .A(\i_iq_demod/demod/QC [0]), .B(
        \i_iq_demod/demod/dp_cluster_0/sub_88/B_not [0]), .Q(
        \i_iq_demod/Q_BB_IN [0]) );
  NAND22 U633 ( .A(\i_iq_demod/filtre_Q/current_state [0]), .B(n1385), .Q(
        \i_iq_demod/filtre_Q/next_state [0]) );
  INV3 U634 ( .A(n1389), .Q(\i_iq_demod/filtre_Q/sel [1]) );
  NAND22 U635 ( .A(n1273), .B(n1268), .Q(
        \i_iq_demod/filtre_Q/out_factor2_req [1]) );
  NAND22 U636 ( .A(n1269), .B(n1270), .Q(
        \i_iq_demod/filtre_Q/out_factor2_req [2]) );
  NOR20 U637 ( .A(n1263), .B(n1264), .Q(n1270) );
  NAND22 U639 ( .A(n1269), .B(n1274), .Q(
        \i_iq_demod/filtre_Q/out_factor2_req [3]) );
  INV0 U640 ( .A(n1264), .Q(n1268) );
  NAND22 U641 ( .A(n1275), .B(n1268), .Q(
        \i_iq_demod/filtre_Q/out_factor1_req [0]) );
  NOR20 U642 ( .A(n1266), .B(n1267), .Q(n1275) );
  NOR31 U643 ( .A(n1266), .B(n1265), .C(n1263), .Q(n289) );
  NAND22 U644 ( .A(n1273), .B(n1274), .Q(
        \i_iq_demod/filtre_Q/out_factor1_req [2]) );
  INV0 U645 ( .A(n1265), .Q(n1273) );
  NAND22 U646 ( .A(n1269), .B(n1274), .Q(
        \i_iq_demod/filtre_Q/out_factor1_req [4]) );
  NAND22 U647 ( .A(n1272), .B(n1274), .Q(
        \i_iq_demod/filtre_Q/out_factor1_req [5]) );
  INV0 U648 ( .A(n1266), .Q(n1272) );
  NAND22 U649 ( .A(n1271), .B(n1274), .Q(
        \i_iq_demod/filtre_Q/out_factor1_req [6]) );
  NOR20 U650 ( .A(n1266), .B(n1267), .Q(n1271) );
  NAND22 U651 ( .A(n1269), .B(n1274), .Q(
        \i_iq_demod/filtre_Q/out_factor1_req [7]) );
  NAND22 U652 ( .A(n1269), .B(n1274), .Q(
        \i_iq_demod/filtre_Q/out_factor1_req [8]) );
  XOR21 U656 ( .A(\i_iq_demod/demod/dp_cluster_1/sub_mult_87/carry [1]), .B(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [1]), .Q(
        \i_iq_demod/I_BB_IN [1]) );
  XOR21 U657 ( .A(\i_iq_demod/demod/IC [0]), .B(\i_iq_demod/demod/QS [0]), .Q(
        \i_iq_demod/I_BB_IN [0]) );
  NAND22 U658 ( .A(\i_iq_demod/filtre_I/current_state [0]), .B(
        \i_iq_demod/filtre_I/n2 ), .Q(\i_iq_demod/filtre_I/next_state [0]) );
  INV3 U659 ( .A(\i_iq_demod/filtre_I/n9 ), .Q(\i_iq_demod/filtre_I/sel [1])
         );
  NAND22 U660 ( .A(\i_iq_demod/filtre_I/factor/n52 ), .B(
        \i_iq_demod/filtre_I/factor/n11 ), .Q(
        \i_iq_demod/filtre_I/out_factor2_req [1]) );
  NAND22 U661 ( .A(\i_iq_demod/filtre_I/factor/n24 ), .B(
        \i_iq_demod/filtre_I/factor/n26 ), .Q(
        \i_iq_demod/filtre_I/out_factor2_req [2]) );
  NOR20 U662 ( .A(\i_iq_demod/filtre_I/factor/n4 ), .B(
        \i_iq_demod/filtre_I/factor/n5 ), .Q(\i_iq_demod/filtre_I/factor/n26 )
         );
  NAND22 U664 ( .A(\i_iq_demod/filtre_I/factor/n24 ), .B(
        \i_iq_demod/filtre_I/factor/n23 ), .Q(
        \i_iq_demod/filtre_I/out_factor2_req [3]) );
  INV0 U665 ( .A(\i_iq_demod/filtre_I/factor/n5 ), .Q(
        \i_iq_demod/filtre_I/factor/n11 ) );
  NAND22 U666 ( .A(\i_iq_demod/filtre_I/factor/n57 ), .B(
        \i_iq_demod/filtre_I/factor/n11 ), .Q(
        \i_iq_demod/filtre_I/out_factor1_req [0]) );
  NOR20 U667 ( .A(\i_iq_demod/filtre_I/factor/n7 ), .B(
        \i_iq_demod/filtre_I/factor/n8 ), .Q(\i_iq_demod/filtre_I/factor/n57 )
         );
  NOR31 U668 ( .A(\i_iq_demod/filtre_I/factor/n7 ), .B(
        \i_iq_demod/filtre_I/factor/n6 ), .C(\i_iq_demod/filtre_I/factor/n4 ), 
        .Q(n290) );
  NAND22 U669 ( .A(\i_iq_demod/filtre_I/factor/n52 ), .B(
        \i_iq_demod/filtre_I/factor/n23 ), .Q(
        \i_iq_demod/filtre_I/out_factor1_req [2]) );
  INV0 U670 ( .A(\i_iq_demod/filtre_I/factor/n6 ), .Q(
        \i_iq_demod/filtre_I/factor/n52 ) );
  NAND22 U671 ( .A(\i_iq_demod/filtre_I/factor/n24 ), .B(
        \i_iq_demod/filtre_I/factor/n23 ), .Q(
        \i_iq_demod/filtre_I/out_factor1_req [4]) );
  NAND22 U672 ( .A(\i_iq_demod/filtre_I/factor/n42 ), .B(
        \i_iq_demod/filtre_I/factor/n23 ), .Q(
        \i_iq_demod/filtre_I/out_factor1_req [5]) );
  INV0 U673 ( .A(\i_iq_demod/filtre_I/factor/n7 ), .Q(
        \i_iq_demod/filtre_I/factor/n42 ) );
  NAND22 U674 ( .A(\i_iq_demod/filtre_I/factor/n39 ), .B(
        \i_iq_demod/filtre_I/factor/n23 ), .Q(
        \i_iq_demod/filtre_I/out_factor1_req [6]) );
  NOR20 U675 ( .A(\i_iq_demod/filtre_I/factor/n7 ), .B(
        \i_iq_demod/filtre_I/factor/n8 ), .Q(\i_iq_demod/filtre_I/factor/n39 )
         );
  NAND22 U676 ( .A(\i_iq_demod/filtre_I/factor/n24 ), .B(
        \i_iq_demod/filtre_I/factor/n23 ), .Q(
        \i_iq_demod/filtre_I/out_factor1_req [7]) );
  NAND22 U677 ( .A(\i_iq_demod/filtre_I/factor/n24 ), .B(
        \i_iq_demod/filtre_I/factor/n23 ), .Q(
        \i_iq_demod/filtre_I/out_factor1_req [8]) );
  NAND22 U678 ( .A(\i_mod_iq/fsm_mapping/n116 ), .B(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/N261 ) );
  NOR31 U679 ( .A(\i_mod_iq/fsm_mapping/n161 ), .B(\i_mod_iq/fsm_mapping/n177 ), .C(\i_mod_iq/fsm_mapping/n166 ), .Q(\i_mod_iq/fsm_mapping/n231 ) );
  NAND22 U680 ( .A(\i_mod_iq/fsm_mapping/n171 ), .B(
        \i_mod_iq/fsm_mapping/N260 ), .Q(\i_mod_iq/fsm_mapping/n168 ) );
  NAND22 U681 ( .A(\i_mod_iq/fsm_mapping/N260 ), .B(
        \i_mod_iq/fsm_mapping/n117 ), .Q(\i_mod_iq/fsm_mapping/n109 ) );
  IMUX40 U682 ( .A(\i_fifo_rx/n533 ), .B(\i_fifo_rx/n523 ), .C(
        \i_fifo_rx/n528 ), .D(\i_fifo_rx/n518 ), .S0(\i_fifo_rx/N44 ), .S1(
        \i_fifo_rx/N43 ), .Q(n291) );
  IMUX40 U683 ( .A(\i_fifo_rx/n513 ), .B(\i_fifo_rx/n503 ), .C(
        \i_fifo_rx/n508 ), .D(\i_fifo_rx/n498 ), .S0(\i_fifo_rx/N44 ), .S1(
        \i_fifo_rx/N43 ), .Q(n292) );
  IMUX40 U684 ( .A(\i_fifo_rx/n493 ), .B(\i_fifo_rx/n483 ), .C(
        \i_fifo_rx/n488 ), .D(\i_fifo_rx/n478 ), .S0(\i_fifo_rx/N44 ), .S1(
        \i_fifo_rx/N43 ), .Q(n293) );
  IMUX40 U685 ( .A(\i_fifo_rx/n473 ), .B(\i_fifo_rx/n463 ), .C(
        \i_fifo_rx/n468 ), .D(\i_fifo_rx/n458 ), .S0(\i_fifo_rx/N44 ), .S1(
        \i_fifo_rx/N43 ), .Q(n294) );
  IMUX40 U686 ( .A(\i_fifo_rx/n453 ), .B(\i_fifo_rx/n443 ), .C(
        \i_fifo_rx/n448 ), .D(\i_fifo_rx/n438 ), .S0(\i_fifo_rx/N44 ), .S1(
        \i_fifo_rx/N43 ), .Q(n295) );
  IMUX40 U687 ( .A(\i_fifo_rx/n433 ), .B(\i_fifo_rx/n423 ), .C(
        \i_fifo_rx/n428 ), .D(\i_fifo_rx/n418 ), .S0(\i_fifo_rx/N44 ), .S1(
        \i_fifo_rx/N43 ), .Q(n296) );
  IMUX40 U688 ( .A(\i_fifo_rx/n413 ), .B(\i_fifo_rx/n403 ), .C(
        \i_fifo_rx/n408 ), .D(\i_fifo_rx/n398 ), .S0(\i_fifo_rx/N44 ), .S1(
        \i_fifo_rx/N43 ), .Q(n297) );
  IMUX40 U689 ( .A(\i_fifo_rx/n393 ), .B(\i_fifo_rx/n383 ), .C(
        \i_fifo_rx/n388 ), .D(\i_fifo_rx/n378 ), .S0(\i_fifo_rx/N44 ), .S1(
        \i_fifo_rx/N43 ), .Q(n298) );
  XOR20 U692 ( .A(\i_fifo_tx/add_180/carry [6]), .B(\i_fifo_tx/rd_ptr[6] ), 
        .Q(\i_fifo_tx/N161 ) );
  XOR20 U693 ( .A(\i_fifo_tx/add_100/carry [6]), .B(\i_fifo_tx/wr_ptr[6] ), 
        .Q(\i_fifo_tx/N134 ) );
  NAND20 U694 ( .A(n317), .B(n126), .Q(n336) );
  NOR20 U695 ( .A(n126), .B(n317), .Q(n337) );
  XNR20 U696 ( .A(\i_fifo_tx/N35 ), .B(\i_fifo_tx/N29 ), .Q(n338) );
  NAND30 U697 ( .A(n340), .B(n339), .C(n338), .Q(n344) );
  XOR20 U698 ( .A(\i_fifo_tx/N34 ), .B(\i_fifo_tx/N28 ), .Q(n343) );
  XOR20 U699 ( .A(\i_fifo_tx/N32 ), .B(\i_fifo_tx/N26 ), .Q(n342) );
  XOR20 U700 ( .A(\i_fifo_tx/N33 ), .B(\i_fifo_tx/N27 ), .Q(n341) );
  NOR40 U701 ( .A(n344), .B(n343), .C(n342), .D(n341), .Q(\i_fifo_tx/N40 ) );
  XOR20 U702 ( .A(\i_fifo_rx/add_139/carry [6]), .B(\i_fifo_rx/rd_ptr[6] ), 
        .Q(\i_fifo_rx/N694 ) );
  XOR20 U703 ( .A(\i_fifo_rx/add_106/carry [6]), .B(\i_fifo_rx/wr_ptr[6] ), 
        .Q(\i_fifo_rx/N86 ) );
  NAND20 U704 ( .A(n302), .B(n133), .Q(n345) );
  NOR20 U705 ( .A(n133), .B(n302), .Q(n346) );
  XNR20 U706 ( .A(\i_fifo_rx/N44 ), .B(\i_fifo_rx/N38 ), .Q(n347) );
  NAND30 U707 ( .A(n349), .B(n348), .C(n347), .Q(n353) );
  XOR20 U708 ( .A(\i_fifo_rx/N43 ), .B(\i_fifo_rx/N37 ), .Q(n352) );
  XOR20 U709 ( .A(\i_fifo_rx/N41 ), .B(\i_fifo_rx/N35 ), .Q(n351) );
  XOR20 U710 ( .A(\i_fifo_rx/N42 ), .B(\i_fifo_rx/N36 ), .Q(n350) );
  NOR40 U711 ( .A(n353), .B(n352), .C(n351), .D(n350), .Q(\i_fifo_rx/N46 ) );
  CLKIN0 U712 ( .A(\i_iq_demod/demod/dp_cluster_1/N85 ), .Q(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [1]) );
  CLKIN0 U713 ( .A(\i_iq_demod/demod/dp_cluster_1/N86 ), .Q(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [2]) );
  CLKIN0 U714 ( .A(\i_iq_demod/demod/dp_cluster_1/N87 ), .Q(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [3]) );
  CLKIN0 U715 ( .A(\i_iq_demod/demod/dp_cluster_1/N88 ), .Q(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [4]) );
  CLKIN0 U716 ( .A(\i_iq_demod/I_BB_IN [0]), .Q(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/carry [1]) );
  CLKIN0 U717 ( .A(\i_iq_demod/demod/dp_cluster_0/N90 ), .Q(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [1]) );
  CLKIN0 U718 ( .A(\i_iq_demod/demod/dp_cluster_0/N91 ), .Q(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [2]) );
  CLKIN0 U719 ( .A(\i_iq_demod/demod/dp_cluster_0/N92 ), .Q(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [3]) );
  CLKIN0 U720 ( .A(\i_iq_demod/demod/dp_cluster_0/N93 ), .Q(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [4]) );
  CLKIN0 U721 ( .A(\i_iq_demod/Q_BB_IN [0]), .Q(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/carry [1]) );
  CLKIN0 U722 ( .A(\i_iq_demod/demod/IS [0]), .Q(
        \i_iq_demod/demod/dp_cluster_0/sub_88/B_not [0]) );
  CLKIN0 U723 ( .A(\i_iq_demod/demod/IS [1]), .Q(
        \i_iq_demod/demod/dp_cluster_0/sub_88/B_not [1]) );
  CLKIN0 U724 ( .A(\i_iq_demod/demod/IS [2]), .Q(
        \i_iq_demod/demod/dp_cluster_0/sub_88/B_not [2]) );
  CLKIN0 U725 ( .A(\i_iq_demod/demod/IS [3]), .Q(
        \i_iq_demod/demod/dp_cluster_0/sub_88/B_not [3]) );
  CLKIN0 U726 ( .A(\i_iq_demod/demod/IS [4]), .Q(
        \i_iq_demod/demod/dp_cluster_0/sub_88/B_not [4]) );
  CLKIN0 U728 ( .A(\i_cordic/cor_y_s0[0][0] ), .Q(
        \i_cordic/S0/sub_50/B_not [0]) );
  CLKIN0 U729 ( .A(\i_cordic/cor_y_s0[0][1] ), .Q(
        \i_cordic/S0/sub_50/B_not [1]) );
  CLKIN0 U730 ( .A(\i_cordic/cor_y_s0[0][2] ), .Q(
        \i_cordic/S0/sub_50/B_not [2]) );
  CLKIN0 U731 ( .A(\i_cordic/cor_y_s0[0][3] ), .Q(
        \i_cordic/S0/sub_50/B_not [3]) );
  CLKIN0 U732 ( .A(\i_cordic/cor_y_s0[0][4] ), .Q(
        \i_cordic/S0/sub_50/B_not [4]) );
  CLKIN0 U733 ( .A(\i_cordic/cor_x_s0[1][2] ), .Q(
        \i_cordic/S1/sub_53/B_not [1]) );
  CLKIN0 U734 ( .A(\i_cordic/cor_x_s0[1][3] ), .Q(
        \i_cordic/S1/sub_53/B_not [2]) );
  CLKIN0 U735 ( .A(\i_cordic/cor_x_s0[1][4] ), .Q(
        \i_cordic/S1/sub_53/B_not [3]) );
  CLKIN0 U736 ( .A(\i_cordic/cor_x_s0[1][5] ), .Q(
        \i_cordic/S1/sub_53/B_not [5]) );
  CLKIN0 U737 ( .A(\i_cordic/cor_y_s0[1][3] ), .Q(
        \i_cordic/S1/sub_50/B_not [2]) );
  CLKIN0 U738 ( .A(\i_cordic/cor_y_s0[1][4] ), .Q(
        \i_cordic/S1/sub_50/B_not [3]) );
  CLKIN0 U739 ( .A(\i_cordic/cor_y_s0[1][1] ), .Q(n354) );
  NOR20 U740 ( .A(n354), .B(\i_cordic/cor_x_s0[1][0] ), .Q(n357) );
  OAI220 U743 ( .A(n357), .B(n360), .C(\i_cordic/cor_y_s0[1][2] ), .D(n356), 
        .Q(\i_cordic/S1/sub_50/carry [2]) );
  CLKIN0 U745 ( .A(\i_cordic/cor_y_s0[1][2] ), .Q(n359) );
  OAI2110 U746 ( .A(\i_cordic/cor_x_s0[1][1] ), .B(\i_cordic/cor_y_s0[1][2] ), 
        .C(\i_cordic/cor_x_s0[1][0] ), .D(\i_cordic/cor_y_s0[1][1] ), .Q(n358)
         );
  OAI210 U747 ( .A(n360), .B(n359), .C(n358), .Q(\i_cordic/S1/add_50/carry [2]) );
  AOI210 U748 ( .A(\i_cordic/cor_y_s1[2][1] ), .B(\i_cordic/cor_x_s1[2][3] ), 
        .C(n361), .Q(n364) );
  CLKIN0 U749 ( .A(n364), .Q(n362) );
  OAI210 U750 ( .A(\i_cordic/cor_y_s1[2][2] ), .B(n362), .C(
        \i_cordic/cor_x_s1[2][4] ), .Q(n363) );
  OAI210 U751 ( .A(n364), .B(n229), .C(n363), .Q(n367) );
  OAI210 U757 ( .A(n370), .B(n236), .C(n369), .Q(\i_cordic/S2/add_53/carry[5] ) );
  NAND20 U758 ( .A(\i_cordic/cor_x_s1[2][2] ), .B(n225), .Q(n372) );
  AOI220 U759 ( .A(n372), .B(\i_cordic/cor_y_s1[2][1] ), .C(n218), .D(n371), 
        .Q(n373) );
  NOR20 U768 ( .A(n260), .B(\i_cdr/i_bit_recovery/phase_q [0]), .Q(n382) );
  OAI220 U769 ( .A(n382), .B(n261), .C(\i_cdr/i_bit_recovery/phase_r [1]), .D(
        n381), .Q(n383) );
  CLKIN0 U770 ( .A(n386), .Q(n384) );
  NOR20 U771 ( .A(\i_cdr/i_bit_recovery/phase_q [3]), .B(n384), .Q(n385) );
  OAI220 U772 ( .A(n386), .B(n262), .C(\i_cdr/i_bit_recovery/phase_r [3]), .D(
        n385), .Q(n387) );
  CLKIN0 U773 ( .A(n387), .Q(n389) );
  NOR20 U774 ( .A(\i_cdr/i_bit_recovery/phase_q [4]), .B(n387), .Q(n388) );
  OAI220 U775 ( .A(n389), .B(n263), .C(\i_cdr/i_bit_recovery/phase_r [4]), .D(
        n388), .Q(\i_cdr/i_bit_recovery/sub_68/carry[5] ) );
  XNR20 U776 ( .A(\i_cdr/i_cdr/cycles[2] ), .B(\i_cdr/i_cdr/count [3]), .Q(
        n393) );
  NOR20 U777 ( .A(\i_cdr/i_cdr/count [1]), .B(n243), .Q(n391) );
  IMUX20 U778 ( .A(n391), .B(n390), .S(\i_cdr/i_cdr/count [2]), .Q(n392) );
  OAI212 U780 ( .A(\i_cdr/i_cdr/n7 ), .B(\i_cdr/i_cdr/n8 ), .C(
        \i_cdr/i_cdr/n9 ), .Q(\i_cdr/i_cdr/n5 ) );
  OAI212 U781 ( .A(\i_iq_demod/gen_sin/current_state [1]), .B(
        \i_iq_demod/gen_sin/current_state [0]), .C(\i_iq_demod/gen_sin/n3 ), 
        .Q(\i_iq_demod/gen_sin/next_state [0]) );
  DFEC3 \i_fifo_rx/rd_ptr_reg[1]  ( .D(\i_fifo_rx/N689 ), .E(\i_fifo_rx/n173 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/N40 ), .QN(n87) );
  ADD31 \i_cordic/S1/add_53/U1_4  ( .A(\i_cordic/cor_y_s0[1][4] ), .B(
        \i_cordic/cor_x_s0[1][5] ), .CI(\i_cordic/S1/add_53/carry [4]), .CO(
        \i_cordic/S1/add_53/carry [5]), .S(\i_cordic/S1/N25 ) );
  XOR31 \i_cordic/S1/sub_50/U2_5  ( .A(\i_cordic/cor_x_s0[1][5] ), .B(
        \i_cordic/S1/sub_50/B_not [5]), .C(\i_cordic/S1/sub_50/carry [5]), .Q(
        \i_cordic/S1/N14 ) );
  DFEC3 \i_fifo_tx/wr_ptr_reg[1]  ( .D(\i_fifo_tx/N129 ), .E(\i_fifo_tx/n152 ), 
        .C(clk_i), .RN(resetn_i), .QN(\i_fifo_tx/n180 ) );
  ADD31 \i_cordic/S1/add_53/U1_3  ( .A(\i_cordic/cor_y_s0[1][3] ), .B(
        \i_cordic/cor_x_s0[1][4] ), .CI(\i_cordic/S1/add_53/carry [3]), .CO(
        \i_cordic/S1/add_53/carry [4]), .S(\i_cordic/S1/N24 ) );
  MUX22 U151 ( .A(n38), .B(n1399), .S(\i_fifo_tx/n153 ), .Q(n1406) );
  IMUX40 U152 ( .A(\i_fifo_tx/n363 ), .B(\i_fifo_tx/n353 ), .C(
        \i_fifo_tx/n358 ), .D(\i_fifo_tx/n348 ), .S0(\i_fifo_tx/N29 ), .S1(
        \i_fifo_tx/N28 ), .Q(n1399) );
  MUX22 U153 ( .A(n39), .B(n1400), .S(\i_fifo_tx/n153 ), .Q(n1408) );
  IMUX40 U154 ( .A(\i_fifo_tx/n343 ), .B(\i_fifo_tx/n333 ), .C(
        \i_fifo_tx/n338 ), .D(\i_fifo_tx/n328 ), .S0(\i_fifo_tx/N29 ), .S1(
        \i_fifo_tx/N28 ), .Q(n1400) );
  MUX22 U155 ( .A(n40), .B(n1401), .S(\i_fifo_tx/n153 ), .Q(n1410) );
  IMUX40 U156 ( .A(\i_fifo_tx/n323 ), .B(\i_fifo_tx/n313 ), .C(
        \i_fifo_tx/n318 ), .D(\i_fifo_tx/n308 ), .S0(\i_fifo_tx/N29 ), .S1(
        \i_fifo_tx/N28 ), .Q(n1401) );
  MUX22 U157 ( .A(n41), .B(n1402), .S(\i_fifo_tx/n153 ), .Q(n1414) );
  IMUX40 U235 ( .A(\i_fifo_tx/n303 ), .B(\i_fifo_tx/n293 ), .C(
        \i_fifo_tx/n298 ), .D(\i_fifo_tx/n288 ), .S0(\i_fifo_tx/N29 ), .S1(
        \i_fifo_tx/N28 ), .Q(n1402) );
  MUX22 U263 ( .A(n42), .B(n1403), .S(\i_fifo_tx/n153 ), .Q(n1418) );
  IMUX40 U264 ( .A(\i_fifo_tx/n283 ), .B(\i_fifo_tx/n273 ), .C(
        \i_fifo_tx/n278 ), .D(\i_fifo_tx/n268 ), .S0(\i_fifo_tx/N29 ), .S1(
        \i_fifo_tx/N28 ), .Q(n1403) );
  MUX22 U266 ( .A(n43), .B(n1404), .S(\i_fifo_tx/n153 ), .Q(n109) );
  IMUX40 U267 ( .A(\i_fifo_tx/n263 ), .B(\i_fifo_tx/n253 ), .C(
        \i_fifo_tx/n258 ), .D(\i_fifo_tx/n248 ), .S0(\i_fifo_tx/N29 ), .S1(
        \i_fifo_tx/N28 ), .Q(n1404) );
  AOI210 U270 ( .A(\i_iq_demod/demod/n32 ), .B(\i_iq_demod/demod/n33 ), .C(
        \i_iq_demod/demod/n31 ), .Q(\i_iq_demod/demod/QC [0]) );
  AOI210 U273 ( .A(\i_iq_demod/demod/n20 ), .B(\i_iq_demod/demod/n22 ), .C(
        \i_iq_demod/demod/n43 ), .Q(\i_iq_demod/demod/IS [0]) );
  NOR21 U274 ( .A(\i_mod_iq/fsm_mapping/n51 ), .B(\i_mod_iq/fsm_mapping/n106 ), 
        .Q(\i_mod_iq/fsm_mapping/n137 ) );
  MUX22 U276 ( .A(\i_iq_demod/filtre_Q/tot [0]), .B(
        \i_iq_demod/filtre_Q/n_temp [0]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N15 ) );
  MUX22 U300 ( .A(\i_iq_demod/filtre_I/tot [0]), .B(
        \i_iq_demod/filtre_I/n_temp [0]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N15 ) );
  XOR31 U301 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[6] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[1][6] ), .C(n968), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][5] ) );
  MUX22 U304 ( .A(\i_iq_demod/filtre_Q/tot [1]), .B(
        \i_iq_demod/filtre_Q/n_temp [1]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N16 ) );
  MUX22 U342 ( .A(\i_iq_demod/filtre_I/tot [1]), .B(
        \i_iq_demod/filtre_I/n_temp [1]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N16 ) );
  XOR31 U344 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[1][6] ), .C(n779), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][5] ) );
  XOR31 U354 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[4] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][4] ), .C(n853), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][3] ) );
  MUX22 U360 ( .A(\i_iq_demod/filtre_Q/tot [2]), .B(
        \i_iq_demod/filtre_Q/n_temp [2]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N17 ) );
  MUX22 U389 ( .A(\i_iq_demod/filtre_I/tot [2]), .B(
        \i_iq_demod/filtre_I/n_temp [2]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N17 ) );
  XOR31 U395 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[6] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][6] ), .C(n1662), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][5] ) );
  MUX22 U452 ( .A(\i_iq_demod/filtre_Q/tot [3]), .B(
        \i_iq_demod/filtre_Q/n_temp [3]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N18 ) );
  MUX22 U460 ( .A(\i_iq_demod/filtre_I/tot [3]), .B(
        \i_iq_demod/filtre_I/n_temp [3]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N18 ) );
  NOR40 U482 ( .A(\i_fifo_rx/n180 ), .B(\i_fifo_rx/n179 ), .C(\i_fifo_rx/n198 ), .D(\i_fifo_rx/n188 ), .Q(\i_fifo_rx/n196 ) );
  XOR31 U484 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[4] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[5] ), .C(n784), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][3] ) );
  XOR31 U489 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_3_net_[4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[5] ), .C(n405), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[2][3] ) );
  XOR31 U491 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][6] ), .C(n870), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[6][5] ) );
  MUX22 U498 ( .A(\i_iq_demod/filtre_Q/tot [4]), .B(
        \i_iq_demod/filtre_Q/n_temp [4]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N19 ) );
  MUX22 U499 ( .A(\i_iq_demod/filtre_I/tot [4]), .B(
        \i_iq_demod/filtre_I/n_temp [4]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N19 ) );
  NOR40 U500 ( .A(\i_fifo_rx/n180 ), .B(\i_fifo_rx/i [0]), .C(\i_fifo_rx/n198 ), .D(\i_fifo_rx/n188 ), .Q(\i_fifo_rx/n194 ) );
  XNR31 U502 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[9] ), .C(n585), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][7] ) );
  XNR31 U505 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[9] ), .C(n396), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[2][7] ) );
  XNR31 U506 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][8] ), .C(n987), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][7] ) );
  XOR31 U541 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][2] ), .C(n693), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[6][1] ) );
  XOR31 U544 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][6] ), .C(n1677), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[6][5] ) );
  IMUX21 U582 ( .A(\i_fifo_rx/shift_register [7]), .B(\i_fifo_rx/N87 ), .S(
        \i_fifo_rx/n170 ), .Q(n1405) );
  XOR31 U584 ( .A(n1232), .B(\i_iq_demod/filtre_Q/tot [6]), .C(
        \i_iq_demod/filtre_Q/temp [6]), .Q(\i_iq_demod/filtre_Q/n_temp [6]) );
  XOR31 U585 ( .A(\i_iq_demod/filtre_I/temp_adder/n7 ), .B(
        \i_iq_demod/filtre_I/tot [6]), .C(\i_iq_demod/filtre_I/temp [6]), .Q(
        \i_iq_demod/filtre_I/n_temp [6]) );
  NOR40 U586 ( .A(\i_fifo_rx/n179 ), .B(\i_fifo_rx/i [1]), .C(\i_fifo_rx/n198 ), .D(\i_fifo_rx/n188 ), .Q(\i_fifo_rx/n192 ) );
  XOR31 U596 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_3_net_[6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[1][6] ), .C(n589), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][5] ) );
  XNR31 U628 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[9] ), .C(n964), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][7] ) );
  XNR31 U630 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_6_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][8] ), .C(n608), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][7] ) );
  XNR31 U653 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][8] ), .C(n1629), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][7] ) );
  XOR31 U763 ( .A(n1178), .B(\i_iq_demod/filtre_Q/mult2 [10]), .C(
        \i_iq_demod/filtre_Q/mult1 [10]), .Q(\i_iq_demod/filtre_Q/tot [10]) );
  XOR31 U764 ( .A(n1171), .B(\i_iq_demod/filtre_Q/mult2 [12]), .C(
        \i_iq_demod/filtre_Q/mult1 [12]), .Q(\i_iq_demod/filtre_Q/tot [12]) );
  XOR31 U765 ( .A(\i_iq_demod/filtre_I/tot_adder/n35 ), .B(
        \i_iq_demod/filtre_I/mult2 [10]), .C(\i_iq_demod/filtre_I/mult1 [10]), 
        .Q(\i_iq_demod/filtre_I/tot [10]) );
  XOR31 U766 ( .A(\i_iq_demod/filtre_I/tot_adder/n28 ), .B(
        \i_iq_demod/filtre_I/mult2 [12]), .C(\i_iq_demod/filtre_I/mult1 [12]), 
        .Q(\i_iq_demod/filtre_I/tot [12]) );
  IMAJ31 U767 ( .A(n376), .B(\i_cordic/cor_y_s1[2][3] ), .C(n226), .Q(n377) );
  IMUX21 U782 ( .A(\i_fifo_rx/shift_register [6]), .B(\i_fifo_rx/N88 ), .S(
        \i_fifo_rx/n170 ), .Q(n1407) );
  XOR31 U784 ( .A(n1228), .B(\i_iq_demod/filtre_Q/tot [8]), .C(
        \i_iq_demod/filtre_Q/temp [8]), .Q(\i_iq_demod/filtre_Q/n_temp [8]) );
  XOR31 U785 ( .A(\i_iq_demod/filtre_I/temp_adder/n3 ), .B(
        \i_iq_demod/filtre_I/tot [8]), .C(\i_iq_demod/filtre_I/temp [8]), .Q(
        \i_iq_demod/filtre_I/n_temp [8]) );
  NOR40 U786 ( .A(\i_fifo_rx/i [0]), .B(\i_fifo_rx/i [1]), .C(\i_fifo_rx/n198 ), .D(\i_fifo_rx/n188 ), .Q(\i_fifo_rx/n189 ) );
  XOR31 U788 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[4] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][4] ), .C(n876), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[6][3] ) );
  XOR31 U793 ( .A(n1086), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[6][4] ), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[4] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[7][3] ) );
  NAND31 U802 ( .A(\i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [2]), .B(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [1]), .C(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/carry [1]), .Q(n102) );
  IMAJ31 U803 ( .A(\i_iq_demod/filtre_Q/mult2 [12]), .B(
        \i_iq_demod/filtre_Q/mult1 [12]), .C(n1171), .Q(n1170) );
  NAND31 U804 ( .A(\i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [2]), .B(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [1]), .C(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/carry [1]), .Q(n103) );
  IMAJ31 U805 ( .A(\i_iq_demod/filtre_I/mult2 [12]), .B(
        \i_iq_demod/filtre_I/mult1 [12]), .C(
        \i_iq_demod/filtre_I/tot_adder/n28 ), .Q(
        \i_iq_demod/filtre_I/tot_adder/n27 ) );
  IMAJ31 U806 ( .A(n367), .B(\i_cordic/cor_y_s1[2][3] ), .C(
        \i_cordic/cor_x_s1[2][5] ), .Q(n370) );
  IMUX21 U807 ( .A(\i_fifo_rx/shift_register [5]), .B(\i_fifo_rx/N89 ), .S(
        \i_fifo_rx/n170 ), .Q(n1409) );
  XOR31 U809 ( .A(n1251), .B(\i_iq_demod/filtre_Q/tot [10]), .C(
        \i_iq_demod/filtre_Q/temp [10]), .Q(\i_iq_demod/filtre_Q/n_temp [10])
         );
  XOR31 U810 ( .A(\i_iq_demod/filtre_I/temp_adder/n42 ), .B(
        \i_iq_demod/filtre_I/tot [10]), .C(\i_iq_demod/filtre_I/temp [10]), 
        .Q(\i_iq_demod/filtre_I/n_temp [10]) );
  NOR40 U811 ( .A(\i_fifo_rx/n179 ), .B(\i_fifo_rx/n180 ), .C(\i_fifo_rx/n188 ), .D(\i_fifo_rx/i [2]), .Q(\i_fifo_rx/n186 ) );
  XOR31 U813 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[4] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][4] ), .C(n830), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][3] ) );
  XOR31 U816 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_21_net_[2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[7][2] ), .C(n727), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[8][1] ) );
  XOR31 U818 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[7][2] ), .B(
        n1625), .C(\i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[2] ), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[8][1] ) );
  XOR31 U820 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[7][2] ), .C(n1106), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[8][1] ) );
  XOR31 U822 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_21_net_[2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[7][2] ), .C(n537), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[8][1] ) );
  NOR21 U825 ( .A(n1411), .B(n1412), .Q(demod_iq_valid_o) );
  NOR31 U826 ( .A(\i_cordic/cor_x_s0[1][1] ), .B(n354), .C(
        \i_cordic/cor_x_s0[1][0] ), .Q(n356) );
  IMUX21 U827 ( .A(\i_fifo_rx/shift_register [4]), .B(\i_fifo_rx/N90 ), .S(
        \i_fifo_rx/n170 ), .Q(n1413) );
  XNR21 U831 ( .A(\i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [4]), .B(
        n119), .Q(\i_iq_demod/Q_BB_IN [4]) );
  MUX22 U832 ( .A(n1389), .B(n1348), .S(\i_iq_demod/filtre_Q/sel [0]), .Q(
        \i_iq_demod/filtre_Q/out_factor2_req [0]) );
  XOR31 U833 ( .A(n1246), .B(\i_iq_demod/filtre_Q/tot [12]), .C(
        \i_iq_demod/filtre_Q/temp [12]), .Q(\i_iq_demod/filtre_Q/n_temp [12])
         );
  XNR21 U834 ( .A(\i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [4]), .B(
        n120), .Q(\i_iq_demod/I_BB_IN [4]) );
  MUX22 U835 ( .A(\i_iq_demod/filtre_I/n9 ), .B(n1311), .S(
        \i_iq_demod/filtre_I/sel [0]), .Q(
        \i_iq_demod/filtre_I/out_factor2_req [0]) );
  XOR31 U836 ( .A(\i_iq_demod/filtre_I/temp_adder/n35 ), .B(
        \i_iq_demod/filtre_I/tot [12]), .C(\i_iq_demod/filtre_I/temp [12]), 
        .Q(\i_iq_demod/filtre_I/n_temp [12]) );
  NOR40 U837 ( .A(\i_fifo_rx/i [0]), .B(\i_fifo_rx/n180 ), .C(\i_fifo_rx/n188 ), .D(\i_fifo_rx/i [2]), .Q(\i_fifo_rx/n184 ) );
  XOR31 U838 ( .A(\i_cordic/cor_y_s1[2][5] ), .B(n226), .C(
        \i_cordic/S2/sub_53/carry[5] ), .Q(\i_cordic/S2/N20 ) );
  XOR31 U841 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[4] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][4] ), .C(n1066), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[6][3] ) );
  XOR31 U846 ( .A(n1166), .B(\i_iq_demod/filtre_Q/mult2 [2]), .C(
        \i_iq_demod/filtre_Q/mult1 [2]), .Q(\i_iq_demod/filtre_Q/tot [2]) );
  XOR31 U847 ( .A(n1162), .B(\i_iq_demod/filtre_Q/mult2 [4]), .C(
        \i_iq_demod/filtre_Q/mult1 [4]), .Q(\i_iq_demod/filtre_Q/tot [4]) );
  XOR31 U848 ( .A(n1158), .B(\i_iq_demod/filtre_Q/mult2 [6]), .C(
        \i_iq_demod/filtre_Q/mult1 [6]), .Q(\i_iq_demod/filtre_Q/tot [6]) );
  XOR31 U849 ( .A(n1154), .B(\i_iq_demod/filtre_Q/mult2 [8]), .C(
        \i_iq_demod/filtre_Q/mult1 [8]), .Q(\i_iq_demod/filtre_Q/tot [8]) );
  XOR31 U850 ( .A(\i_iq_demod/filtre_I/tot_adder/n15 ), .B(
        \i_iq_demod/filtre_I/mult2 [2]), .C(\i_iq_demod/filtre_I/mult1 [2]), 
        .Q(\i_iq_demod/filtre_I/tot [2]) );
  XOR31 U851 ( .A(\i_iq_demod/filtre_I/tot_adder/n11 ), .B(
        \i_iq_demod/filtre_I/mult2 [4]), .C(\i_iq_demod/filtre_I/mult1 [4]), 
        .Q(\i_iq_demod/filtre_I/tot [4]) );
  XOR31 U852 ( .A(\i_iq_demod/filtre_I/tot_adder/n7 ), .B(
        \i_iq_demod/filtre_I/mult2 [6]), .C(\i_iq_demod/filtre_I/mult1 [6]), 
        .Q(\i_iq_demod/filtre_I/tot [6]) );
  XOR31 U853 ( .A(\i_iq_demod/filtre_I/tot_adder/n3 ), .B(
        \i_iq_demod/filtre_I/mult2 [8]), .C(\i_iq_demod/filtre_I/mult1 [8]), 
        .Q(\i_iq_demod/filtre_I/tot [8]) );
  IMUX21 U854 ( .A(\i_fifo_rx/shift_register [3]), .B(\i_fifo_rx/N91 ), .S(
        \i_fifo_rx/n170 ), .Q(n1417) );
  XOR31 U858 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[8][2] ), .B(
        n1665), .C(\i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[2] ), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[9][1] ) );
  XOR31 U859 ( .A(n1663), .B(n1738), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[2] ), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[9][1] ) );
  XNR21 U860 ( .A(n102), .B(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [3]), .Q(
        \i_iq_demod/Q_BB_IN [3]) );
  XNR21 U861 ( .A(n110), .B(
        \i_iq_demod/demod/dp_cluster_0/sub_mult_88/B_not [2]), .Q(
        \i_iq_demod/Q_BB_IN [2]) );
  MUX22 U863 ( .A(\i_iq_demod/filtre_Q/tot [13]), .B(
        \i_iq_demod/filtre_Q/n_temp [13]), .S(n1391), .Q(
        \i_iq_demod/filtre_Q/N28 ) );
  XOR31 U865 ( .A(n550), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[8][2] ), .C(
        \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[2] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[9][1] ) );
  XNR21 U866 ( .A(n103), .B(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [3]), .Q(
        \i_iq_demod/I_BB_IN [3]) );
  XNR21 U867 ( .A(n111), .B(
        \i_iq_demod/demod/dp_cluster_1/sub_mult_87/B_not [2]), .Q(
        \i_iq_demod/I_BB_IN [2]) );
  MUX22 U869 ( .A(\i_iq_demod/filtre_I/tot [13]), .B(
        \i_iq_demod/filtre_I/n_temp [13]), .S(\i_iq_demod/filtre_I/n22 ), .Q(
        \i_iq_demod/filtre_I/N28 ) );
  NOR40 U870 ( .A(\i_fifo_rx/i [1]), .B(\i_fifo_rx/n179 ), .C(\i_fifo_rx/n188 ), .D(\i_fifo_rx/i [2]), .Q(\i_fifo_rx/n182 ) );
  XOR21 U872 ( .A(\i_cordic/S2/N31 ), .B(n329), .Q(\i_cordic/S2/N37 ) );
  OAI222 U874 ( .A(n499), .B(n500), .C(n501), .D(n502), .Q(n497) );
  OAI222 U875 ( .A(n547), .B(n500), .C(n549), .D(n548), .Q(n544) );
  OAI222 U886 ( .A(n832), .B(n833), .C(n834), .D(n1935), .Q(n830) );
  OAI222 U888 ( .A(n1543), .B(n856), .C(n857), .D(n1932), .Q(n853) );
  OAI222 U889 ( .A(n786), .B(n787), .C(n789), .D(n788), .Q(n784) );
  OAI222 U904 ( .A(n596), .B(n597), .C(n599), .D(n598), .Q(n594) );
  NOR31 U907 ( .A(\i_iq_demod/filtre_I/sel [0]), .B(
        \i_iq_demod/filtre_I/sel [1]), .C(n1311), .Q(
        \i_iq_demod/filtre_I/data_reg1/n7 ) );
  NOR31 U908 ( .A(\i_iq_demod/filtre_Q/sel [0]), .B(
        \i_iq_demod/filtre_Q/sel [1]), .C(n1348), .Q(n1318) );
  NOR31 U909 ( .A(\i_iq_demod/filtre_I/sel [0]), .B(
        \i_iq_demod/filtre_I/sel [1]), .C(n1311), .Q(n1282) );
  NOR31 U910 ( .A(\i_iq_demod/filtre_Q/sel [0]), .B(
        \i_iq_demod/filtre_Q/sel [1]), .C(n1348), .Q(n1355) );
  NOR31 U913 ( .A(\i_iq_demod/filtre_I/sel [1]), .B(
        \i_iq_demod/filtre_I/sel [2]), .C(\i_iq_demod/filtre_I/data_reg1/n36 ), 
        .Q(\i_iq_demod/filtre_I/data_reg1/n4 ) );
  NOR31 U914 ( .A(\i_iq_demod/filtre_Q/sel [1]), .B(
        \i_iq_demod/filtre_Q/sel [2]), .C(n1347), .Q(n1315) );
  NOR31 U916 ( .A(\i_iq_demod/filtre_I/sel [1]), .B(n1943), .C(
        \i_iq_demod/filtre_I/data_reg1/n36 ), .Q(n1279) );
  NOR31 U917 ( .A(\i_iq_demod/filtre_Q/sel [1]), .B(n1944), .C(n1347), .Q(
        n1352) );
  OAI221 U923 ( .A(N10), .B(n36), .C(n47), .D(n191), .Q(fifo_rx_data_i) );
  NAND22 U926 ( .A(\i_iq_demod/cosine_IN [0]), .B(\i_iq_demod/gen_sin/n3 ), 
        .Q(\i_iq_demod/demod/n33 ) );
  INV3 U930 ( .A(\i_mod_iq/fsm_mapping/n65 ), .Q(\i_mod_iq/fsm_mapping/n194 )
         );
  NAND22 U931 ( .A(\i_mod_iq/fsm_mapping/n188 ), .B(\i_mod_iq/fsm_mapping/n69 ), .Q(\i_mod_iq/fsm_mapping/n187 ) );
  IMUX21 U932 ( .A(\i_cordic/S2/n37 ), .B(\i_cordic/S2/n37 ), .S(
        \i_cordic/S2/n21 ), .Q(\i_cordic/cor_w_s1[4][2] ) );
  INV3 U933 ( .A(\i_cordic/S2/n36 ), .Q(\i_cordic/S3/N36 ) );
  IMUX21 U934 ( .A(\i_cordic/S2/n34 ), .B(\i_cordic/S2/n34 ), .S(
        \i_cordic/S2/n21 ), .Q(\i_cordic/cor_w_s1[4][5] ) );
  DFEC3 \i_fifo_tx/rd_ptr_reg[0]  ( .D(n126), .E(\i_fifo_tx/n187 ), .C(clk_i), 
        .RN(resetn_i), .Q(\i_fifo_tx/N30 ), .QN(n126) );
  DFEC3 \i_fifo_rx/rd_ptr_reg[0]  ( .D(n133), .E(\i_fifo_rx/n173 ), .C(clk_i), 
        .RN(resetn_i), .Q(\i_fifo_rx/N39 ), .QN(n133) );
  DFEC3 \i_fifo_tx/rd_ptr_reg[3]  ( .D(\i_fifo_tx/N158 ), .E(\i_fifo_tx/n187 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/N33 ), .QN(n269) );
  DFEC3 \i_fifo_rx/rd_ptr_reg[3]  ( .D(\i_fifo_rx/N691 ), .E(\i_fifo_rx/n173 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/N42 ), .QN(n271) );
  DFEC1 \i_fifo_tx/wr_ptr_reg[2]  ( .D(\i_fifo_tx/N130 ), .E(\i_fifo_tx/n152 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/N26 ), .QN(\i_fifo_tx/n182 )
         );
  ADD21 \i_fifo_tx/add_100/U1_1_2  ( .A(n1946), .B(
        \i_fifo_tx/add_100/carry [2]), .CO(\i_fifo_tx/add_100/carry [3]), .S(
        \i_fifo_tx/N130 ) );
  DFEC1 \i_fifo_rx/wr_ptr_reg[2]  ( .D(\i_fifo_rx/N82 ), .E(\i_fifo_rx/n171 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/N35 ), .QN(\i_fifo_rx/n155 )
         );
  ADD21 \i_fifo_rx/add_106/U1_1_2  ( .A(n1945), .B(
        \i_fifo_rx/add_106/carry [2]), .CO(\i_fifo_rx/add_106/carry [3]), .S(
        \i_fifo_rx/N82 ) );
  DFC3 \i_cordic/ibb_ibuff_reg[4]  ( .D(cordic_ibb_i[4]), .C(clk_i), .RN(
        resetn_i), .Q(\i_cordic/S0/N32 ), .QN(\i_cordic/n5 ) );
  DFEC1 \i_fifo_tx/rd_ptr_reg[2]  ( .D(\i_fifo_tx/N157 ), .E(\i_fifo_tx/n187 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/N32 ), .QN(n1940) );
  ADD21 \i_fifo_tx/add_180/U1_1_2  ( .A(n1941), .B(
        \i_fifo_tx/add_180/carry [2]), .CO(\i_fifo_tx/add_180/carry [3]), .S(
        \i_fifo_tx/N157 ) );
  DFEC1 \i_fifo_rx/rd_ptr_reg[2]  ( .D(\i_fifo_rx/N690 ), .E(\i_fifo_rx/n173 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/N41 ), .QN(n1938) );
  XOR31 \i_cordic/S2/add_53/U1_5  ( .A(\i_cordic/cor_y_s1[2][5] ), .B(
        \i_cordic/cor_x_s1[2][5] ), .C(\i_cordic/S2/add_53/carry[5] ), .Q(
        \i_cordic/S2/N26 ) );
  DFEC3 \i_fifo_rx/wr_ptr_reg[0]  ( .D(\i_fifo_rx/n154 ), .E(\i_fifo_rx/n171 ), 
        .C(clk_i), .RN(resetn_i), .Q(n134), .QN(\i_fifo_rx/n154 ) );
  DFEC3 \i_fifo_tx/wr_ptr_reg[0]  ( .D(\i_fifo_tx/n181 ), .E(\i_fifo_tx/n152 ), 
        .C(clk_i), .RN(resetn_i), .Q(n132), .QN(\i_fifo_tx/n181 ) );
  DFEC3 \i_fifo_tx/rd_ptr_reg[5]  ( .D(\i_fifo_tx/N160 ), .E(\i_fifo_tx/n187 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/N35 ) );
  DFEC3 \i_fifo_rx/wr_ptr_reg[4]  ( .D(\i_fifo_rx/N84 ), .E(\i_fifo_rx/n171 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/N37 ), .QN(\i_fifo_rx/n45 ) );
  DFEC3 \i_fifo_tx/wr_ptr_reg[4]  ( .D(\i_fifo_tx/N132 ), .E(\i_fifo_tx/n152 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/N28 ), .QN(\i_fifo_tx/n170 )
         );
  DFEC3 \i_fifo_rx/rd_ptr_reg[5]  ( .D(\i_fifo_rx/N693 ), .E(\i_fifo_rx/n173 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/N44 ) );
  DFEC3 \i_fifo_rx/wr_ptr_reg[1]  ( .D(\i_fifo_rx/N81 ), .E(\i_fifo_rx/n171 ), 
        .C(clk_i), .RN(resetn_i), .Q(n86), .QN(\i_fifo_rx/n153 ) );
  DFEC3 \i_fifo_rx/wr_ptr_reg[3]  ( .D(\i_fifo_rx/N83 ), .E(\i_fifo_rx/n171 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_rx/N36 ), .QN(\i_fifo_rx/n46 ) );
  DFEC3 \i_fifo_tx/wr_ptr_reg[3]  ( .D(\i_fifo_tx/N131 ), .E(\i_fifo_tx/n152 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/N27 ), .QN(\i_fifo_tx/n171 )
         );
  DFEC3 \i_fifo_tx/rd_ptr_reg[4]  ( .D(\i_fifo_tx/N159 ), .E(\i_fifo_tx/n187 ), 
        .C(clk_i), .RN(resetn_i), .Q(\i_fifo_tx/N34 ) );
  ADD21 \i_fifo_rx/add_139/U1_1_4  ( .A(\i_fifo_rx/N43 ), .B(
        \i_fifo_rx/add_139/carry [4]), .CO(\i_fifo_rx/add_139/carry [5]), .S(
        \i_fifo_rx/N692 ) );
  DFC3 \i_iq_demod/filtre_I/data_1_1_reg[0]  ( .D(
        \i_iq_demod/filtre_I/data_1_1_req [0]), .C(clk_i), .RN(resetn_i), .Q(
        net41341), .QN(n164) );
  DFC3 \i_iq_demod/filtre_Q/data_1_1_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/data_1_1_req [0]), .C(clk_i), .RN(resetn_i), .Q(
        n1920), .QN(n162) );
  DFC3 \i_iq_demod/filtre_Q/out_factor1_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1_req [2]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_Q/out_factor1 [2]), .QN(n199) );
  DFC3 \i_iq_demod/filtre_I/out_factor1_reg[1]  ( .D(
        \i_iq_demod/filtre_I/out_factor1_req [1]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_I/out_factor1 [1]), .QN(n202) );
  DFC3 \i_iq_demod/filtre_Q/data_2_1_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/data_2_1_req [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_2_1 [1]), .QN(n1917) );
  DFC3 \i_iq_demod/filtre_Q/data_1_1_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/data_1_1_req [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_1_1 [1]), .QN(n1916) );
  DFC3 \i_iq_demod/filtre_I/data_2_1_reg[1]  ( .D(
        \i_iq_demod/filtre_I/data_2_1_req [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_2_1 [1]), .QN(n1924) );
  DFC3 \i_iq_demod/filtre_I/data_1_1_reg[1]  ( .D(
        \i_iq_demod/filtre_I/data_1_1_req [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_1_1 [1]), .QN(n1923) );
  DFC3 \i_iq_demod/filtre_I/out_factor1_reg[2]  ( .D(
        \i_iq_demod/filtre_I/out_factor1_req [2]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_I/out_factor1 [2]), .QN(n201) );
  DFC3 \i_iq_demod/filtre_I/data_2_1_reg[0]  ( .D(
        \i_iq_demod/filtre_I/data_2_1_req [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_2_1 [0]), .QN(n198) );
  DFC3 \i_iq_demod/filtre_I/data_1_2_reg[0]  ( .D(
        \i_iq_demod/filtre_I/data_1_2_req [0]), .C(clk_i), .RN(resetn_i), .Q(
        n1882), .QN(n161) );
  DFC3 \i_iq_demod/filtre_Q/data_1_2_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/data_1_2_req [0]), .C(clk_i), .RN(resetn_i), .Q(
        n1861), .QN(n163) );
  DFC3 \i_iq_demod/filtre_Q/out_factor1_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1_req [1]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_Q/out_factor1 [1]), .QN(n200) );
  DFC3 \i_iq_demod/filtre_Q/data_2_1_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/data_2_1_req [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_2_1 [0]), .QN(n196) );
  DFC3 \i_iq_demod/filtre_I/data_2_2_reg[1]  ( .D(
        \i_iq_demod/filtre_I/data_2_2_req [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_2_2 [1]), .QN(n1873) );
  DFC3 \i_iq_demod/filtre_I/data_1_2_reg[1]  ( .D(
        \i_iq_demod/filtre_I/data_1_2_req [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_1_2 [1]), .QN(n1524) );
  DFC3 \i_iq_demod/filtre_Q/out_factor2_reg[2]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2_req [2]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_Q/out_factor2 [2]), .QN(n152) );
  DFC3 \i_iq_demod/filtre_Q/data_2_2_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/data_2_2_req [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_2_2 [1]) );
  DFC3 \i_iq_demod/filtre_I/out_factor2_reg[2]  ( .D(
        \i_iq_demod/filtre_I/out_factor2_req [2]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_I/out_factor2 [2]), .QN(n148) );
  DFC3 \i_iq_demod/filtre_Q/data_1_2_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/data_1_2_req [1]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_1_2 [1]) );
  DFC3 \i_iq_demod/filtre_I/out_factor1_reg[4]  ( .D(
        \i_iq_demod/filtre_I/out_factor1_req [4]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_I/out_factor1 [4]), .QN(n154) );
  DFC3 \i_iq_demod/filtre_I/out_factor2_reg[1]  ( .D(
        \i_iq_demod/filtre_I/out_factor2_req [1]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_I/out_factor2 [1]), .QN(n149) );
  DFC3 \i_iq_demod/filtre_I/out_factor1_reg[3]  ( .D(
        \i_iq_demod/filtre_I/out_factor1_req [3]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_I/out_factor1 [3]), .QN(n130) );
  DFC3 \i_iq_demod/filtre_I/data_2_2_reg[0]  ( .D(
        \i_iq_demod/filtre_I/data_2_2_req [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_I/data_2_2 [0]), .QN(n195) );
  DFC3 \i_iq_demod/filtre_Q/data_2_2_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/data_2_2_req [0]), .C(clk_i), .RN(resetn_i), .Q(
        \i_iq_demod/filtre_Q/data_2_2 [0]), .QN(n197) );
  DFC3 \i_iq_demod/filtre_Q/out_factor2_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2_req [3]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_Q/out_factor2 [3]), .QN(n128) );
  DFC3 \i_iq_demod/filtre_Q/out_factor1_reg[3]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1_req [3]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_Q/out_factor1 [3]), .QN(n127) );
  DFC3 \i_iq_demod/filtre_Q/out_factor2_reg[1]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2_req [1]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_Q/out_factor2 [1]), .QN(n153) );
  DFC3 \i_iq_demod/filtre_Q/out_factor2_reg[0]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2_req [0]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_Q/out_factor2 [0]), .QN(n145) );
  DFC3 \i_iq_demod/filtre_I/out_factor2_reg[3]  ( .D(
        \i_iq_demod/filtre_I/out_factor2_req [3]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_I/out_factor2 [3]), .QN(n131) );
  DFC3 \i_iq_demod/filtre_I/out_factor2_reg[4]  ( .D(
        \i_iq_demod/filtre_I/out_factor2_req [4]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_I/out_factor2 [4]), .QN(n147) );
  DFC3 \i_iq_demod/filtre_Q/out_factor2_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/out_factor2_req [4]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_Q/out_factor2 [4]), .QN(n151) );
  DFC3 \i_iq_demod/filtre_Q/out_factor1_reg[4]  ( .D(
        \i_iq_demod/filtre_Q/out_factor1_req [4]), .C(clk_i), .RN(resetn_i), 
        .Q(\i_iq_demod/filtre_Q/out_factor1 [4]), .QN(n150) );
  XOR31 U753 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_18_net_[4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[6][4] ), .C(n517), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[7][3] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U96  ( .A(n130), .B(n174), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[3] ) );
  XOR31 U798 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_21_net_[4] ), .B(n532), .C(n1455), .Q(\i_iq_demod/filtre_I/mult1_multiplier/register[8][3] ) );
  NOR20 \i_iq_demod/filtre_I/mult1_multiplier/U64  ( .A(n142), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[5] ) );
  XNR20 \i_iq_demod/filtre_I/mult1_multiplier/genblk1[2].adder/U39  ( .A(n439), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/register[2][0] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/S_pipe [2]) );
  OAI222 U879 ( .A(n431), .B(n432), .C(net41468), .D(n433), .Q(n429) );
  IMAJ31 U245 ( .A(n1592), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[2] ), .C(n435), .Q(n433)
         );
  DFEC3 \i_mod_iq/fsm_mapping/cpt_reg[2]  ( .D(\i_mod_iq/fsm_mapping/n37 ), 
        .E(\i_mod_iq/fsm_mapping/n183 ), .C(clk_i), .RN(resetn_i), .Q(
        \i_mod_iq/fsm_mapping/cpt [2]), .QN(\i_mod_iq/fsm_mapping/n69 ) );
  NAND24 U162 ( .A(n1822), .B(n1823), .Q(n711) );
  BUF6 U163 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][2] ), .Q(
        n1419) );
  BUF6 U164 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_0_net_[3] ), .Q(n1664)
         );
  INV6 U165 ( .A(n1675), .Q(n1676) );
  NOR24 U170 ( .A(n201), .B(n1829), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[2] ) );
  NAND23 U171 ( .A(\i_iq_demod/filtre_I/data_2_2 [1]), .B(
        \i_iq_demod/filtre_I/data_1_2 [1]), .Q(n1878) );
  CLKIN6 U172 ( .A(n1071), .Q(n1497) );
  INV4 U173 ( .A(n1579), .Q(n529) );
  BUF15 U174 ( .A(n1416), .Q(n1615) );
  BUF6 U175 ( .A(n645), .Q(n1420) );
  NOR21 U176 ( .A(n128), .B(n1771), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[3] ) );
  NAND24 U177 ( .A(n1870), .B(n1871), .Q(n536) );
  XOR22 U178 ( .A(net41707), .B(n1588), .Q(n1455) );
  NAND24 U179 ( .A(n1495), .B(n1496), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[6][4] ) );
  CLKIN6 U186 ( .A(n1888), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][3] ) );
  MAJ32 U189 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[4][6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[6] ), .C(n658), .Q(
        n1694) );
  XOR22 U190 ( .A(n1674), .B(n1487), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][1] ) );
  XNR22 U191 ( .A(n990), .B(n989), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][6] ) );
  NAND26 U193 ( .A(n1796), .B(n1797), .Q(n1025) );
  INV6 U194 ( .A(n1429), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][1] ) );
  NAND26 U195 ( .A(n1803), .B(n1802), .Q(n1869) );
  NOR22 U196 ( .A(n507), .B(n524), .Q(n527) );
  NOR22 U197 ( .A(n127), .B(n1729), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[3] ) );
  NAND20 U199 ( .A(n1745), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[1] ), .Q(n1009) );
  XOR22 U200 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[3] ), .Q(n1487) );
  NAND21 U205 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][3] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[3] ), .Q(n1872) );
  CLKIN6 U208 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][3] ), .Q(
        n1600) );
  CLKIN6 U210 ( .A(n1858), .Q(n927) );
  CLKBU15 U211 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[6][4] ), 
        .Q(n1518) );
  NAND22 U212 ( .A(n1523), .B(n497), .Q(n1469) );
  CLKIN3 U216 ( .A(n997), .Q(n1754) );
  AOI222 U217 ( .A(n1722), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[7] ), .C(n1710), .D(n823), .Q(n821) );
  XOR22 U218 ( .A(n828), .B(n1913), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][4] ) );
  XNR22 U219 ( .A(n874), .B(n1928), .Q(n1608) );
  BUF8 U220 ( .A(n875), .Q(n1928) );
  CLKIN12 U221 ( .A(n1645), .Q(n896) );
  MAJ32 U222 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[3][6] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[6] ), .C(n446), .Q(
        net42883) );
  CLKIN6 U234 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[6][5] ), .Q(
        n1883) );
  AOI221 U237 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_15_net_[7] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[5][7] ), .C(n1435), .D(
        n489), .Q(n487) );
  NAND24 U240 ( .A(n1808), .B(n1809), .Q(n549) );
  NOR23 U242 ( .A(n149), .B(n135), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[1] ) );
  CLKIN4 U244 ( .A(n1784), .Q(n135) );
  NAND34 U247 ( .A(net42278), .B(net42279), .C(n1445), .Q(n1572) );
  MAJ32 U249 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[6][4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[4] ), .C(n517), .Q(
        n1445) );
  BUF4 U250 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][4] ), .Q(
        n1707) );
  NAND24 U255 ( .A(n1464), .B(n1465), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[6][4] ) );
  CLKIN2 U256 ( .A(n1445), .Q(n1588) );
  NAND21 U269 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[8][3] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[3] ), .Q(n1808) );
  CLKIN1 U271 ( .A(n977), .Q(n1509) );
  NOR22 U272 ( .A(n130), .B(n1709), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[3] ) );
  NAND24 U279 ( .A(n1225), .B(n1223), .Q(n1488) );
  MAJ32 U280 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][6] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[6] ), .C(n468), .Q(
        net42758) );
  NAND33 U283 ( .A(n1416), .B(\i_iq_demod/filtre_Q/out_factor2 [1]), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[2] ), .Q(n1884) );
  XOR22 U287 ( .A(n1862), .B(\i_iq_demod/filtre_Q/data_2_2 [0]), .Q(n137) );
  CLKIN6 U303 ( .A(n1861), .Q(n1862) );
  MAJ32 U306 ( .A(n1518), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[4] ), .C(n707), .Q(
        n1649) );
  NOR24 U307 ( .A(n152), .B(n137), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[2] ) );
  XNR22 U308 ( .A(n1753), .B(n1702), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][5] ) );
  CLKIN6 U310 ( .A(n825), .Q(n1702) );
  XOR22 U312 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][6] ), .Q(n1753) );
  XNR22 U314 ( .A(n824), .B(n823), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][6] ) );
  INV6 U317 ( .A(n1520), .Q(n1749) );
  INV0 U318 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[3][0] ), .Q(
        n838) );
  NAND24 U319 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[3][0] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[0] ), .Q(n1480) );
  XNR22 U320 ( .A(n1893), .B(n820), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][0] ) );
  XNR22 U325 ( .A(n1531), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[4] ), .Q(n1044) );
  XNR22 U326 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][1] ), .Q(n1075) );
  INV6 U328 ( .A(n1705), .Q(n1084) );
  MAJ32 U330 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[6][4] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[4] ), .C(n1086), .Q(
        n1705) );
  XOR22 U334 ( .A(n1812), .B(n1857), .Q(n1727) );
  BUF8 U335 ( .A(n995), .Q(n1812) );
  XNR22 U348 ( .A(n1528), .B(n1033), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][7] ) );
  AOI222 U350 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[4][7] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[7] ), .C(n1733), .D(
        n1035), .Q(n1033) );
  NAND26 U351 ( .A(n1787), .B(n1110), .Q(n1106) );
  XNR22 U352 ( .A(n1649), .B(n706), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[7][4] ) );
  XNR22 U355 ( .A(n684), .B(n1883), .Q(n706) );
  NAND24 U358 ( .A(n1875), .B(n1876), .Q(n1911) );
  XOR22 U361 ( .A(n1921), .B(\i_iq_demod/filtre_Q/data_2_1 [0]), .Q(n1728) );
  CLKIN6 U364 ( .A(n1920), .Q(n1921) );
  CLKIN6 U365 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[5][5] ), .Q(
        n1540) );
  CLKIN4 U367 ( .A(n1612), .Q(n1653) );
  XOR22 U369 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[7][4] ), .B(
        n1616), .Q(n1612) );
  XNR22 U375 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_0_net_[4] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[3] ), .Q(n599) );
  AOI222 U378 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[7] ), .C(n1725), .D(n777), .Q(n775) );
  MAJ32 U382 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[1][6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[6] ), .C(n779), .Q(n1725) );
  XOR22 U384 ( .A(n1749), .B(n1869), .Q(n1531) );
  INV4 U385 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[3] ), .Q(n1506)
         );
  NAND24 U386 ( .A(n1505), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[3] ), .Q(n1508) );
  NOR22 U392 ( .A(n128), .B(n1671), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[3] ) );
  NOR21 U400 ( .A(n151), .B(n1671), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[4] ) );
  NAND26 U403 ( .A(n1503), .B(n1504), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][4] ) );
  CLKBU12 U406 ( .A(n1830), .Q(n1857) );
  BUF6 U410 ( .A(n204), .Q(n1671) );
  NAND24 U411 ( .A(n1795), .B(n1799), .Q(n1797) );
  NAND22 U412 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][5] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[5] ), .Q(n1886) );
  NAND24 U414 ( .A(n1908), .B(net41535), .Q(net41468) );
  INV3 U415 ( .A(n1713), .Q(n616) );
  INV3 U416 ( .A(n1800), .Q(n639) );
  XOR21 U417 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[6] ), .Q(n1491) );
  XOR21 U418 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[6] ), .Q(n1466) );
  BUF8 U421 ( .A(n1636), .Q(n1892) );
  NAND22 U422 ( .A(n1552), .B(n1857), .Q(n1555) );
  INV3 U423 ( .A(n1812), .Q(n1552) );
  NAND23 U424 ( .A(n1756), .B(n1757), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][3] ) );
  NAND22 U425 ( .A(n1754), .B(n1755), .Q(n1757) );
  NOR21 U429 ( .A(n151), .B(n1770), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[4] ) );
  BUF2 U437 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[2][4] ), .Q(
        n1606) );
  INV3 U438 ( .A(n1827), .Q(n635) );
  NAND23 U439 ( .A(n1543), .B(n856), .Q(n1545) );
  XNR21 U441 ( .A(n1044), .B(n1043), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][3] ) );
  NAND24 U443 ( .A(n1507), .B(n1508), .Q(n1003) );
  XOR21 U446 ( .A(n1699), .B(n1013), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][6] ) );
  NAND26 U447 ( .A(n1872), .B(net41833), .Q(net41781) );
  NOR21 U449 ( .A(n156), .B(\i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[6] ) );
  NAND24 U454 ( .A(n1470), .B(n1471), .Q(n1582) );
  NAND22 U457 ( .A(n1724), .B(n667), .Q(n1876) );
  AOI221 U459 ( .A(n1696), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[7] ), .C(n1827), .D(n634), .Q(n632) );
  NAND22 U461 ( .A(n1563), .B(n690), .Q(n1823) );
  INV3 U469 ( .A(n857), .Q(n1667) );
  INV3 U470 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][0] ), .Q(
        n816) );
  INV3 U471 ( .A(n1786), .Q(n880) );
  XOR21 U472 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][3] ), .B(
        n1866), .Q(n1071) );
  INV3 U473 ( .A(n1457), .Q(n1731) );
  INV3 U479 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[1] ), .Q(n1763)
         );
  NOR22 U481 ( .A(n152), .B(n1774), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[2] ) );
  NAND22 U483 ( .A(n1538), .B(n1539), .Q(n1090) );
  NAND22 U485 ( .A(n1701), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[3] ), .Q(n1538) );
  INV3 U487 ( .A(net41468), .Q(net43481) );
  NOR22 U490 ( .A(n130), .B(n138), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[3] ) );
  INV3 U492 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_15_net_[6] ), .Q(n1587) );
  NAND22 U494 ( .A(n1567), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[5] ), .Q(net42278) );
  XOR21 U501 ( .A(n1582), .B(n1583), .Q(n1567) );
  NAND22 U503 ( .A(net42278), .B(net42279), .Q(net41707) );
  NAND33 U504 ( .A(n1513), .B(n1514), .C(n1515), .Q(n1516) );
  INV3 U507 ( .A(n697), .Q(n1515) );
  XOR21 U509 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[5][7] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[7] ), .Q(n679) );
  NOR23 U511 ( .A(n199), .B(n1728), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[2] ) );
  MAJ31 U512 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[5][6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[6] ), .C(n870), .Q(
        n1609) );
  NOR21 U513 ( .A(n150), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[4] ) );
  NAND22 U514 ( .A(n1615), .B(\i_iq_demod/filtre_Q/out_factor2 [2]), .Q(n1643)
         );
  BUF2 U515 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[3] ), .Q(n1638)
         );
  XOR21 U517 ( .A(n1089), .B(n1670), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[7][2] ) );
  NAND22 U519 ( .A(n1567), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[5] ), .Q(n1571) );
  INV3 U520 ( .A(net41341), .Q(n1590) );
  CLKIN3 U521 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_0_net_[1] ), .Q(n602) );
  INV3 U527 ( .A(n722), .Q(n1842) );
  NOR21 U528 ( .A(n143), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[0] ) );
  NAND22 U529 ( .A(n1816), .B(n1929), .Q(n1818) );
  NAND23 U530 ( .A(n1838), .B(n1895), .Q(n1839) );
  INV3 U531 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[1] ), .Q(n1895)
         );
  INV3 U532 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][1] ), .Q(
        n1838) );
  XNR21 U533 ( .A(n1216), .B(n1214), .Q(n1915) );
  NAND22 U534 ( .A(n1678), .B(n1926), .Q(n1860) );
  NAND22 U545 ( .A(n1859), .B(n1860), .Q(n1906) );
  INV3 U546 ( .A(n1721), .Q(n899) );
  NAND24 U547 ( .A(n1550), .B(n1551), .Q(n1052) );
  XOR21 U548 ( .A(n1853), .B(n1010), .Q(n1718) );
  NOR21 U549 ( .A(n128), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[3] ) );
  NAND22 U550 ( .A(n1764), .B(net42565), .Q(n438) );
  INV3 U573 ( .A(n1584), .Q(n1576) );
  NAND23 U574 ( .A(n534), .B(n1930), .Q(n1871) );
  INV6 U575 ( .A(\i_fifo_tx/n171 ), .Q(n273) );
  INV6 U576 ( .A(\i_fifo_rx/n46 ), .Q(n274) );
  NAND24 U577 ( .A(\i_iq_demod/filtre_I/out_factor2 [0]), .B(n1716), .Q(n1715)
         );
  NAND24 U578 ( .A(n1844), .B(n1843), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[8][3] ) );
  NAND22 U579 ( .A(n1842), .B(n1653), .Q(n1844) );
  NAND22 U580 ( .A(n722), .B(n1612), .Q(n1843) );
  NAND23 U581 ( .A(n1840), .B(n1841), .Q(n1845) );
  NAND23 U583 ( .A(n908), .B(n1926), .Q(n1841) );
  BUF2 U589 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[8][2] ), .Q(
        n1663) );
  NAND22 U590 ( .A(n1475), .B(n1476), .Q(n1477) );
  INV3 U592 ( .A(\i_iq_demod/filtre_I/_15_net_[8] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/n25 ) );
  XNR21 U593 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[8][4] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[4] ), .Q(n736) );
  OAI222 U594 ( .A(n1620), .B(n1637), .C(n995), .D(n1830), .Q(n1662) );
  BUF2 U595 ( .A(n993), .Q(n1620) );
  XOR21 U597 ( .A(n1725), .B(n777), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][6] ) );
  MAJ32 U614 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[4][5] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[5] ), .C(n1863), .Q(
        n658) );
  MUX24 U617 ( .A(net42078), .B(net43270), .S(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[3] ), .Q(n1898) );
  NOR23 U621 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][6] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[6] ), .Q(n1421) );
  INV6 U623 ( .A(n1421), .Q(n1471) );
  NAND23 U625 ( .A(n1557), .B(n1852), .Q(n1559) );
  OAI312 U629 ( .A(n482), .B(n484), .C(n483), .D(n485), .Q(n480) );
  MUX21 U638 ( .A(\i_cordic/S0/r64/carry [5]), .B(\i_cordic/S0/N14 ), .S(n1942), .Q(\i_cordic/cor_x_s0[1][5] ) );
  OAI222 U654 ( .A(n975), .B(n1837), .C(n978), .D(n977), .Q(n973) );
  INV3 U655 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[4] ), .Q(n975)
         );
  OAI222 U663 ( .A(n804), .B(n805), .C(n806), .D(n807), .Q(n802) );
  INV3 U690 ( .A(n1889), .Q(n806) );
  NOR21 U691 ( .A(n1671), .B(n141), .Q(n1422) );
  INV3 U727 ( .A(n1422), .Q(n1637) );
  NOR21 U741 ( .A(n166), .B(n130), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[3] ) );
  MAJ31 U742 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][3] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[3] ), .C(n1654), .Q(
        n1066) );
  XOR22 U744 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][5] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[5] ), .Q(net41996) );
  NAND22 U752 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][0] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[0] ), .Q(n1423) );
  INV3 U754 ( .A(n1423), .Q(n1500) );
  OAI222 U755 ( .A(n683), .B(n684), .C(n685), .D(n686), .Q(n1677) );
  INV3 U756 ( .A(n1630), .Q(n685) );
  NAND31 U760 ( .A(\i_iq_demod/filtre_I/out_factor1 [1]), .B(n1424), .C(
        \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[2] ), .Q(n416) );
  INV3 U761 ( .A(n1709), .Q(n1424) );
  XNR31 U762 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_9_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][8] ), .C(n442), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][7] ) );
  XNR22 U779 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][2] ), .Q(n1027) );
  OAI222 U783 ( .A(n1564), .B(n879), .C(n914), .D(n915), .Q(n911) );
  CLKIN6 U787 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[7][3] ), .Q(
        n1564) );
  OAI222 U789 ( .A(\i_cordic/S0/n39 ), .B(n277), .C(
        \i_cordic/S0/sub_53/carry [5]), .D(n1942), .Q(
        \i_cordic/cor_y_s0[1][5] ) );
  NOR21 U790 ( .A(n1766), .B(n141), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[5] ) );
  INV3 U791 ( .A(n1615), .Q(n1766) );
  XNR31 U792 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[9] ), .C(n775), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][7] ) );
  OAI222 U794 ( .A(n1865), .B(n1805), .C(n1047), .D(n1864), .Q(n1043) );
  INV3 U795 ( .A(n1644), .Q(n1047) );
  XNR21 U796 ( .A(n1863), .B(n663), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][4] ) );
  MAJ32 U797 ( .A(n1419), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[2] ), .C(n859), .Q(
        n1425) );
  INV3 U799 ( .A(n1425), .Q(n857) );
  NAND21 U800 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[1] ), .Q(n630) );
  OAI311 U801 ( .A(n714), .B(n697), .C(n715), .D(n716), .Q(n712) );
  OAI212 U808 ( .A(n1075), .B(n1499), .C(n1077), .Q(n1072) );
  XOR21 U812 ( .A(n1609), .B(n868), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[6][6] ) );
  OAI312 U814 ( .A(n413), .B(n415), .C(n414), .D(n416), .Q(n1934) );
  CLKIN3 U815 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_3_net_[0] ), .Q(n415) );
  CLKIN6 U817 ( .A(net41344), .Q(n414) );
  NAND22 U819 ( .A(n1583), .B(n1580), .Q(n1574) );
  INV2 U821 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][6] ), .Q(
        n1580) );
  INV3 U823 ( .A(n1719), .Q(n914) );
  XOR22 U824 ( .A(n1004), .B(n1896), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][1] ) );
  NOR21 U828 ( .A(n174), .B(n146), .Q(n1426) );
  INV3 U829 ( .A(n1426), .Q(n484) );
  MUX21 U830 ( .A(\i_cordic/S1/N8 ), .B(\i_cordic/S1/N14 ), .S(
        \i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/cor_x_s0[2][5] ) );
  XNR21 U839 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][5] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[5] ), .Q(n617) );
  OAI212 U840 ( .A(n1467), .B(n1692), .C(n1468), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][6] ) );
  INV3 U842 ( .A(n800), .Q(n1467) );
  NOR21 U843 ( .A(n1766), .B(n176), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[9] ) );
  XOR31 U844 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_6_net_[4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[2][4] ), .C(n429), .Q(
        n1427) );
  INV3 U845 ( .A(n1427), .Q(net42078) );
  XNR22 U855 ( .A(n1603), .B(n1599), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[5][4] ) );
  XOR21 U856 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[4] ), .B(n1632), .Q(n1428) );
  INV3 U857 ( .A(n1428), .Q(n789) );
  NOR21 U862 ( .A(n152), .B(n210), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[2] ) );
  NAND22 U864 ( .A(n1569), .B(n1589), .Q(net42279) );
  NAND24 U868 ( .A(n1516), .B(n698), .Q(n693) );
  XNR31 U871 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_3_net_[2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[3] ), .C(n1912), .Q(
        n1429) );
  XNR21 U873 ( .A(n686), .B(n1630), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[6][4] ) );
  XNR22 U876 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][2] ), .Q(n883) );
  NOR23 U877 ( .A(n1890), .B(n200), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[1] ) );
  NAND21 U878 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[7][1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[1] ), .Q(n1110) );
  CLKIN3 U880 ( .A(n1439), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[7][1] ) );
  INV3 U881 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_0_net_[1] ), .Q(n413)
         );
  MAJ31 U882 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[6][6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[6] ), .C(n890), .Q(
        n1769) );
  XNR21 U883 ( .A(n1220), .B(n1219), .Q(n1430) );
  INV3 U884 ( .A(n1430), .Q(n206) );
  MUX21 U885 ( .A(\i_cordic/S1/N7 ), .B(\i_cordic/S1/N13 ), .S(
        \i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/cor_x_s0[2][4] ) );
  NOR20 U887 ( .A(n193), .B(n169), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[6] ) );
  CLKIN6 U890 ( .A(n1415), .Q(n193) );
  XNR22 U891 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[4] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][4] ), .Q(n999) );
  NAND22 U892 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][0] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[0] ), .Q(n1499) );
  XNR31 U893 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_9_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][8] ), .C(n632), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][7] ) );
  XNR21 U894 ( .A(n1863), .B(n663), .Q(n1685) );
  NAND22 U895 ( .A(n1915), .B(\i_iq_demod/filtre_Q/out_factor1 [2]), .Q(n1431)
         );
  INV3 U896 ( .A(n1431), .Q(\i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[2] )
         );
  OAI212 U897 ( .A(n1608), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[4] ), .C(n1556), .Q(
        n1619) );
  MAJ32 U898 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[6][2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[2] ), .C(n1091), .Q(
        n1432) );
  INV3 U899 ( .A(n1432), .Q(n1089) );
  NAND21 U900 ( .A(net41398), .B(net41996), .Q(n1464) );
  OAI312 U901 ( .A(n1433), .B(n1434), .C(n730), .D(n731), .Q(n727) );
  INV3 U902 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[7][0] ), .Q(
        n1433) );
  INV3 U903 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[0] ), .Q(n1434) );
  NAND22 U905 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[2][1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[1] ), .Q(net42565) );
  INV3 U906 ( .A(n1933), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[2][1] ) );
  XOR22 U911 ( .A(n1581), .B(n1584), .Q(n1586) );
  XNR22 U912 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[6][1] ), .Q(n904) );
  INV3 U915 ( .A(n1573), .Q(n1435) );
  NOR21 U918 ( .A(n651), .B(n1634), .Q(n653) );
  XNR31 U919 ( .A(n1769), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[6][7] ), .C(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[7] ), .Q(n1910) );
  XNR20 U920 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[1] ), .Q(n1607) );
  NAND22 U921 ( .A(\i_iq_demod/filtre_I/out_factor1 [0]), .B(n1443), .Q(n461)
         );
  XNR30 U922 ( .A(\i_cordic/cor_y_s0[1][5] ), .B(\i_cordic/cor_x_s0[1][5] ), 
        .C(\i_cordic/S1/sub_53/carry [5]), .Q(\i_cordic/S1/N20 ) );
  NAND22 U924 ( .A(n1502), .B(n972), .Q(n1503) );
  XOR31 U925 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_3_net_[6] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[1][6] ), .C(n400), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[2][5] ) );
  XOR21 U927 ( .A(n782), .B(n783), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][4] ) );
  NOR21 U928 ( .A(n170), .B(n204), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[6] ) );
  NAND24 U929 ( .A(n1866), .B(n1537), .Q(n1539) );
  INV6 U935 ( .A(n1701), .Q(n1537) );
  XOR30 U936 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[6] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][6] ), .C(n1037), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][5] ) );
  XNR22 U937 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_15_net_[4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[5][4] ), .Q(n1523) );
  XNR31 U938 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][8] ), .C(n821), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][7] ) );
  NAND22 U939 ( .A(n1784), .B(\i_iq_demod/filtre_I/out_factor2 [2]), .Q(n1436)
         );
  INV3 U940 ( .A(n1436), .Q(\i_iq_demod/filtre_I/mult2_multiplier/_0_net_[2] )
         );
  XOR31 U941 ( .A(\i_iq_demod/filtre_I/data_1_2 [2]), .B(
        \i_iq_demod/filtre_I/data_2_2 [2]), .C(n1203), .Q(n1437) );
  INV3 U942 ( .A(n1437), .Q(n203) );
  OAI212 U943 ( .A(n1916), .B(n1917), .C(n1463), .Q(n1212) );
  OAI212 U944 ( .A(n1225), .B(n1223), .C(n1488), .Q(n1416) );
  NOR21 U945 ( .A(n168), .B(n202), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[1] ) );
  XNR21 U946 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_3_net_[2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[3] ), .Q(n1562) );
  NAND22 U947 ( .A(n1817), .B(n1818), .Q(n862) );
  XOR31 U948 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[4] ), .B(
        n1536), .C(n1906), .Q(n1438) );
  INV3 U949 ( .A(n1438), .Q(n1902) );
  XNR31 U950 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[6][2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[2] ), .C(n1091), .Q(
        n1439) );
  NAND22 U951 ( .A(n1549), .B(n1732), .Q(n1551) );
  XOR31 U952 ( .A(\i_iq_demod/filtre_I/sum1_adder/n4 ), .B(
        \i_iq_demod/filtre_I/data_2_1 [4]), .C(
        \i_iq_demod/filtre_I/data_1_1 [4]), .Q(n174) );
  NAND30 U953 ( .A(n1572), .B(n1584), .C(n1571), .Q(n1577) );
  NAND22 U954 ( .A(\i_iq_demod/filtre_I/out_factor2 [0]), .B(n1451), .Q(n674)
         );
  XOR22 U955 ( .A(n909), .B(n1845), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[8][4] ) );
  NAND22 U956 ( .A(\i_iq_demod/filtre_I/out_factor1 [0]), .B(n1593), .Q(n439)
         );
  MUX22 U957 ( .A(\i_cordic/S0/N4 ), .B(\i_cordic/S0/N10 ), .S(
        \i_cordic/cor_y_s0[0][5] ), .Q(\i_cordic/cor_x_s0[1][1] ) );
  MUX21 U958 ( .A(\i_cordic/S1/N20 ), .B(\i_cordic/S1/N26 ), .S(
        \i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/cor_y_s0[2][5] ) );
  MAJ32 U959 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][5] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[5] ), .C(n1713), .Q(n612) );
  NOR22 U960 ( .A(n193), .B(n131), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[3] ) );
  XOR22 U961 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[4] ), .B(n1837), .Q(n978) );
  XNR21 U962 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_0_net_[4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[3] ), .Q(n410) );
  INV3 U963 ( .A(net42230), .Q(net41398) );
  OAI222 U964 ( .A(n690), .B(n1712), .C(n710), .D(n711), .Q(n707) );
  INV3 U965 ( .A(n1706), .Q(n710) );
  XOR31 U966 ( .A(\i_iq_demod/filtre_Q/data_1_1 [2]), .B(
        \i_iq_demod/filtre_Q/data_2_1 [2]), .C(n1212), .Q(n1440) );
  INV3 U967 ( .A(n1440), .Q(n1890) );
  OAI212 U968 ( .A(n1695), .B(n1497), .C(n1498), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[6][2] ) );
  NAND20 U969 ( .A(\i_iq_demod/filtre_Q/data_1_2 [1]), .B(
        \i_iq_demod/filtre_Q/data_2_2 [1]), .Q(n1224) );
  XNR21 U970 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[7][1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[1] ), .Q(n730) );
  NAND23 U971 ( .A(n1776), .B(n1775), .Q(n1777) );
  XNR21 U972 ( .A(n1920), .B(\i_iq_demod/filtre_Q/data_2_1 [0]), .Q(n136) );
  AOI212 U973 ( .A(n1416), .B(\i_iq_demod/filtre_Q/out_factor2 [1]), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[2] ), .Q(n1441) );
  INV3 U974 ( .A(n1441), .Q(n1885) );
  XOR31 U975 ( .A(n1804), .B(n1058), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[6] ), .Q(n1442) );
  INV3 U976 ( .A(n1442), .Q(n1082) );
  OAI212 U977 ( .A(n202), .B(n166), .C(n1933), .Q(n1764) );
  XNR21 U978 ( .A(\i_iq_demod/filtre_I/sum1_adder/n7 ), .B(
        \i_iq_demod/filtre_I/sum1_adder/n6 ), .Q(n1443) );
  INV3 U979 ( .A(n1443), .Q(n168) );
  XNR21 U980 ( .A(n603), .B(n606), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][0] ) );
  XOR21 U981 ( .A(n1719), .B(n1927), .Q(n1444) );
  INV3 U982 ( .A(n1444), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[8][2] ) );
  NOR21 U983 ( .A(n1030), .B(n1718), .Q(n1032) );
  NOR31 U984 ( .A(\i_iq_demod/filtre_I/sel [1]), .B(n1311), .C(
        \i_iq_demod/filtre_I/sel [0]), .Q(\i_iq_demod/filtre_I/factor/n7 ) );
  INV2 U985 ( .A(\i_iq_demod/filtre_I/sel [2]), .Q(n1311) );
  OAI220 U986 ( .A(n909), .B(n1845), .C(n908), .D(n873), .Q(n907) );
  INV3 U987 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[7][5] ), .Q(
        n908) );
  XOR20 U988 ( .A(\i_cordic/cor_y_s0[1][0] ), .B(\i_cordic/cor_x_s0[1][1] ), 
        .Q(\i_cordic/S1/N21 ) );
  XOR21 U989 ( .A(n612), .B(n1466), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][5] ) );
  NOR21 U990 ( .A(n151), .B(n210), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[4] ) );
  XNR22 U991 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[3][3] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[3] ), .Q(n646) );
  XOR31 U992 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[6] ), .C(n847), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][5] ) );
  XNR31 U993 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_6_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[2][8] ), .C(n419), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][7] ) );
  NAND24 U994 ( .A(n1806), .B(n1807), .Q(n686) );
  XNR21 U995 ( .A(n1644), .B(n1864), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][2] ) );
  NOR21 U996 ( .A(n168), .B(n201), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[2] ) );
  NAND22 U997 ( .A(n1207), .B(n1205), .Q(n1824) );
  INV3 U998 ( .A(n1881), .Q(n1207) );
  XNR31 U999 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_12_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][8] ), .C(n654), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][7] ) );
  OAI212 U1000 ( .A(n1560), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][2] ), .C(n1561), .Q(
        n1896) );
  OAI222 U1001 ( .A(n1866), .B(n1735), .C(n1105), .D(n1104), .Q(n1101) );
  NAND22 U1002 ( .A(n1532), .B(\i_iq_demod/filtre_I/_15_net_[8] ), .Q(n1581)
         );
  NOR21 U1003 ( .A(n697), .B(n714), .Q(n717) );
  XNR21 U1004 ( .A(n1521), .B(n631), .Q(n1634) );
  NAND21 U1005 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[0] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][0] ), .Q(n1446) );
  INV3 U1006 ( .A(n1446), .Q(n820) );
  XNR21 U1007 ( .A(n1920), .B(\i_iq_demod/filtre_Q/data_2_1 [0]), .Q(n1729) );
  XOR31 U1008 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[7][1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[1] ), .C(n1111), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[8][0] ) );
  XOR20 U1009 ( .A(n1745), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[1] ), .Q(n1447) );
  INV3 U1010 ( .A(n1447), .Q(n1853) );
  XOR21 U1011 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[7][5] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[5] ), .Q(n1448) );
  INV3 U1012 ( .A(n1448), .Q(n1100) );
  NOR21 U1013 ( .A(n439), .B(n437), .Q(n441) );
  IMUX21 U1014 ( .A(\i_mod_iq/fsm_mapping/n140 ), .B(
        \i_mod_iq/fsm_mapping/n139 ), .S(\i_mod_iq/fsm_mapping/n80 ), .Q(
        \i_mod_iq/fsm_mapping/n135 ) );
  NOR20 U1015 ( .A(n135), .B(n143), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[0] ) );
  XOR31 U1016 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[6] ), .B(
        n1910), .C(n907), .Q(n1618) );
  XOR31 U1017 ( .A(n1240), .B(\i_iq_demod/filtre_Q/tot [2]), .C(
        \i_iq_demod/filtre_Q/temp [2]), .Q(\i_iq_demod/filtre_Q/n_temp [2]) );
  NOR20 U1018 ( .A(n138), .B(n146), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[0] ) );
  CLKIN6 U1019 ( .A(n1826), .Q(n138) );
  XOR31 U1020 ( .A(\i_iq_demod/filtre_I/temp_adder/n15 ), .B(
        \i_iq_demod/filtre_I/tot [2]), .C(\i_iq_demod/filtre_I/temp [2]), .Q(
        \i_iq_demod/filtre_I/n_temp [2]) );
  IMUX21 U1021 ( .A(\i_cordic/n5 ), .B(\i_cordic/S0/N32 ), .S(
        \i_cordic/cor_y_s0[0][5] ), .Q(\i_cordic/S1/N38 ) );
  XNR21 U1022 ( .A(n1657), .B(n398), .Q(n1675) );
  MAJ32 U1023 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[3][5] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[5] ), .C(n1800), .Q(n636) );
  XNR21 U1024 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][7] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[7] ), .Q(n1449) );
  INV3 U1025 ( .A(n1449), .Q(n845) );
  OAI212 U1026 ( .A(n1523), .B(n497), .C(n1469), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[6][3] ) );
  NAND22 U1027 ( .A(n496), .B(net42230), .Q(n1465) );
  NAND33 U1028 ( .A(n1878), .B(n1879), .C(n1881), .Q(n1825) );
  XNR21 U1029 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[6][2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[2] ), .Q(n902) );
  OAI222 U1030 ( .A(n1063), .B(n1525), .C(n1084), .D(n1085), .Q(n1080) );
  NOR21 U1031 ( .A(n1923), .B(n1924), .Q(n1450) );
  INV3 U1032 ( .A(n1450), .Q(\i_iq_demod/filtre_I/sum1_adder/n14 ) );
  XNR31 U1033 ( .A(n1199), .B(\i_iq_demod/filtre_I/data_2_2 [4]), .C(
        \i_iq_demod/filtre_I/data_1_2 [4]), .Q(n1451) );
  INV3 U1034 ( .A(n1451), .Q(n209) );
  XOR20 U1035 ( .A(n1649), .B(n706), .Q(n1648) );
  NAND22 U1036 ( .A(n1565), .B(n1566), .Q(n1927) );
  NOR21 U1037 ( .A(\i_iq_demod/filtre_Q/current_state [1]), .B(
        \i_iq_demod/filtre_Q/current_state [0]), .Q(n1384) );
  NOR21 U1038 ( .A(\i_iq_demod/filtre_I/current_state [1]), .B(
        \i_iq_demod/filtre_I/current_state [0]), .Q(\i_iq_demod/filtre_I/n1 )
         );
  XOR21 U1039 ( .A(n726), .B(n725), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[8][2] ) );
  NOR21 U1040 ( .A(n863), .B(n861), .Q(n865) );
  INV3 U1041 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[0] ), .Q(n863) );
  NOR21 U1042 ( .A(n792), .B(n1658), .Q(n796) );
  INV3 U1043 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[1] ), .Q(n792)
         );
  NOR21 U1044 ( .A(n1076), .B(n1093), .Q(n1096) );
  INV3 U1045 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[6][0] ), .Q(
        n1093) );
  NAND22 U1046 ( .A(\i_iq_demod/filtre_Q/out_factor2 [0]), .B(n1452), .Q(n1008) );
  INV3 U1047 ( .A(n1774), .Q(n1452) );
  XNR21 U1048 ( .A(n1861), .B(\i_iq_demod/filtre_Q/data_2_2 [0]), .Q(n1770) );
  NAND24 U1049 ( .A(n1484), .B(n1485), .Q(n1118) );
  XNR20 U1050 ( .A(n483), .B(n486), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[5][0] ) );
  OAI212 U1051 ( .A(n1475), .B(n1476), .C(n1477), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[2][0] ) );
  AOI221 U1052 ( .A(n1576), .B(n1570), .C(n1578), .D(n1577), .Q(n510) );
  INV3 U1053 ( .A(n1581), .Q(n1578) );
  OAI311 U1054 ( .A(\i_cordic/cor_y_s1[2][4] ), .B(n367), .C(
        \i_cordic/cor_y_s1[2][3] ), .D(\i_cordic/cor_x_s1[2][5] ), .Q(n369) );
  XNR21 U1055 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_9_net_[0] ), .B(
        n1634), .Q(\i_iq_demod/filtre_I/mult2_multiplier/S_pipe [3]) );
  NOR21 U1056 ( .A(n697), .B(n742), .Q(n745) );
  INV3 U1057 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[0] ), .Q(n697) );
  XOR31 U1058 ( .A(n1236), .B(\i_iq_demod/filtre_Q/tot [4]), .C(
        \i_iq_demod/filtre_Q/temp [4]), .Q(\i_iq_demod/filtre_Q/n_temp [4]) );
  XOR31 U1059 ( .A(\i_iq_demod/filtre_I/temp_adder/n11 ), .B(
        \i_iq_demod/filtre_I/tot [4]), .C(\i_iq_demod/filtre_I/temp [4]), .Q(
        \i_iq_demod/filtre_I/n_temp [4]) );
  IMUX20 U1060 ( .A(\i_mod_iq/fsm_mapping/temp_IBB [3]), .B(
        \i_mod_iq/fsm_mapping/n48 ), .S(\i_mod_iq/fsm_mapping/n58 ), .Q(
        \i_mod_iq/fsm_mapping/n50 ) );
  MAJ31 U1061 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[5][6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[6] ), .C(n1677), .Q(
        n1453) );
  XOR21 U1062 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_12_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][8] ), .Q(n1454) );
  NOR21 U1063 ( .A(n147), .B(n135), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[4] ) );
  NOR21 U1064 ( .A(n154), .B(n1709), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[4] ) );
  AOI221 U1065 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[4][7] ), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/_12_net_[7] ), .C(n1694), .D(
        n656), .Q(n654) );
  XNR21 U1066 ( .A(n715), .B(n717), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[7][0] ) );
  CLKIN6 U1067 ( .A(n1603), .Q(n472) );
  NAND26 U1068 ( .A(n1473), .B(n1474), .Q(n1584) );
  XOR21 U1069 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][7] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[7] ), .Q(n489) );
  INV3 U1070 ( .A(n489), .Q(n1472) );
  INV3 U1071 ( .A(n1737), .Q(n1041) );
  INV6 U1072 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][3] ), .Q(
        n1795) );
  INV3 U1073 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[2][3] ), .Q(
        n431) );
  INV6 U1074 ( .A(n1760), .Q(n1761) );
  INV3 U1075 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_6_net_[0] ), .Q(n629)
         );
  XOR21 U1076 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_9_net_[4] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][4] ), .Q(n1456) );
  INV3 U1077 ( .A(n1654), .Q(n1695) );
  INV3 U1078 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][0] ), .Q(
        n1074) );
  IMAJ31 U1079 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][2] ), 
        .B(n1660), .C(n1026), .Q(n1457) );
  NAND22 U1080 ( .A(n1602), .B(n444), .Q(n1460) );
  NAND23 U1081 ( .A(n1458), .B(n1459), .Q(n1461) );
  NAND24 U1082 ( .A(n1460), .B(n1461), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][6] ) );
  CLKIN3 U1083 ( .A(n1602), .Q(n1458) );
  INV3 U1084 ( .A(n444), .Q(n1459) );
  NAND31 U1085 ( .A(n1462), .B(\i_iq_demod/filtre_Q/data_2_1 [0]), .C(n1920), 
        .Q(n1463) );
  INV3 U1086 ( .A(n1214), .Q(n1462) );
  CLKIN6 U1087 ( .A(net41996), .Q(n496) );
  NAND22 U1088 ( .A(n1467), .B(n1692), .Q(n1468) );
  AOI222 U1089 ( .A(n1621), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[7] ), .C(net42883), .D(
        n444), .Q(n442) );
  XNR22 U1090 ( .A(n1456), .B(n1720), .Q(n1724) );
  BUF6 U1091 ( .A(n641), .Q(n1720) );
  INV3 U1092 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[6][3] ), .Q(
        n1848) );
  AOI221 U1093 ( .A(\i_iq_demod/filtre_I/data_2_1 [3]), .B(
        \i_iq_demod/filtre_I/data_1_1 [3]), .C(
        \i_iq_demod/filtre_I/sum1_adder/n5 ), .D(
        \i_iq_demod/filtre_I/sum1_adder/n6 ), .Q(
        \i_iq_demod/filtre_I/sum1_adder/n4 ) );
  XNR21 U1094 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[5] ), .Q(n783) );
  NAND22 U1095 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][6] ), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/_15_net_[6] ), .Q(n1470) );
  NAND22 U1096 ( .A(n489), .B(n1585), .Q(n1473) );
  NAND26 U1097 ( .A(n1472), .B(n1573), .Q(n1474) );
  INV3 U1098 ( .A(net41786), .Q(n1475) );
  INV3 U1099 ( .A(n417), .Q(n1476) );
  XOR21 U1100 ( .A(n1919), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[6] ), .Q(n1478) );
  XOR21 U1101 ( .A(n1097), .B(n1478), .Q(n1821) );
  OAI220 U1102 ( .A(n1098), .B(n1063), .C(n1517), .D(n1100), .Q(n1097) );
  NOR21 U1103 ( .A(n149), .B(n203), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[1] ) );
  XOR22 U1104 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][6] ), .B(
        n1698), .Q(n1479) );
  XOR22 U1105 ( .A(n1814), .B(n1479), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[6][5] ) );
  NAND23 U1106 ( .A(n1522), .B(n1481), .Q(n1903) );
  INV3 U1107 ( .A(n1480), .Q(n1481) );
  NAND23 U1108 ( .A(n1903), .B(n841), .Q(n836) );
  NAND22 U1109 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[8][3] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[3] ), .Q(n1484) );
  NAND28 U1110 ( .A(n1482), .B(n1483), .Q(n1485) );
  CLKIN6 U1111 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[8][3] ), 
        .Q(n1482) );
  INV15 U1112 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[3] ), .Q(
        n1483) );
  XOR21 U1113 ( .A(\i_iq_demod/filtre_Q/data_1_2 [2]), .B(n1611), .Q(n1486) );
  XOR21 U1114 ( .A(n1767), .B(n1486), .Q(n1641) );
  NOR21 U1115 ( .A(n153), .B(n1641), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[1] ) );
  NOR22 U1116 ( .A(n163), .B(n197), .Q(n1225) );
  XOR21 U1117 ( .A(\i_iq_demod/filtre_I/data_1_1 [2]), .B(
        \i_iq_demod/filtre_I/data_2_1 [2]), .Q(n1489) );
  XOR22 U1118 ( .A(n1596), .B(n1489), .Q(n1593) );
  INV6 U1119 ( .A(n1593), .Q(n166) );
  XOR22 U1120 ( .A(n1638), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[2] ), .Q(n1490) );
  XOR22 U1121 ( .A(n979), .B(n1490), .Q(n1745) );
  INV3 U1122 ( .A(n1643), .Q(\i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[2] ) );
  OAI311 U1123 ( .A(n981), .B(n1772), .C(n982), .D(n1884), .Q(n979) );
  XOR22 U1124 ( .A(n802), .B(n1491), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][5] ) );
  NOR21 U1125 ( .A(n150), .B(n136), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[4] ) );
  XNR22 U1126 ( .A(n1454), .B(n464), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[5][7] ) );
  XOR22 U1127 ( .A(n1639), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[4] ), .Q(n1492) );
  XOR22 U1128 ( .A(n1020), .B(n1492), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][3] ) );
  NAND21 U1129 ( .A(n1907), .B(n1494), .Q(n1495) );
  NAND22 U1130 ( .A(n1493), .B(n1064), .Q(n1496) );
  CLKIN1 U1131 ( .A(n1907), .Q(n1493) );
  INV1 U1132 ( .A(n1064), .Q(n1494) );
  NAND22 U1133 ( .A(n1695), .B(n1497), .Q(n1498) );
  NAND24 U1134 ( .A(n1521), .B(n1500), .Q(n1880) );
  NAND22 U1135 ( .A(n1501), .B(n1686), .Q(n1504) );
  CLKIN1 U1136 ( .A(n972), .Q(n1501) );
  CLKIN6 U1137 ( .A(n1686), .Q(n1502) );
  NAND22 U1138 ( .A(n1900), .B(n1506), .Q(n1507) );
  CLKIN3 U1139 ( .A(n1900), .Q(n1505) );
  NAND20 U1140 ( .A(n977), .B(n1510), .Q(n1511) );
  NAND22 U1141 ( .A(n1509), .B(n978), .Q(n1512) );
  NAND22 U1142 ( .A(n1511), .B(n1512), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][2] ) );
  INV2 U1143 ( .A(n978), .Q(n1510) );
  CLKBU6 U1144 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[2][2] ), 
        .Q(n1744) );
  NAND22 U1145 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[2][2] ), 
        .B(n1560), .Q(n1561) );
  CLKIN3 U1146 ( .A(n695), .Q(n1513) );
  CLKIN6 U1147 ( .A(n696), .Q(n1514) );
  CLKIN3 U1148 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[5][0] ), 
        .Q(n695) );
  NAND21 U1149 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][1] ), .Q(n698) );
  MAJ32 U1150 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[5][2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[2] ), .C(n693), .Q(
        n1768) );
  NAND26 U1151 ( .A(n1880), .B(n630), .Q(n625) );
  CLKIN1 U1152 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[8][3] ), 
        .Q(n737) );
  OAI311 U1153 ( .A(n1052), .B(n1051), .C(n1053), .D(n1054), .Q(n1739) );
  XNR20 U1154 ( .A(n673), .B(n676), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][0] ) );
  XNR20 U1155 ( .A(n1113), .B(n1115), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[9][3] ) );
  NAND22 U1156 ( .A(n1690), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[3] ), .Q(n1822) );
  XNR22 U1157 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[8][4] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[4] ), .Q(n1115) );
  XOR22 U1158 ( .A(n1517), .B(n1100), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[8][4] ) );
  CLKIN6 U1159 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][5] ), 
        .Q(n1016) );
  CLKIN6 U1160 ( .A(n1060), .Q(n1814) );
  NAND23 U1161 ( .A(n1882), .B(\i_iq_demod/filtre_I/data_2_2 [0]), .Q(n1881)
         );
  BUF6 U1162 ( .A(n1530), .Q(n1517) );
  MAJ32 U1163 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][6] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[6] ), .C(n1060), .Q(
        n1804) );
  XNR30 U1164 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[6] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][6] ), .C(n1060), .Q(
        n1525) );
  NAND24 U1165 ( .A(n1887), .B(n1886), .Q(n1907) );
  XNR20 U1166 ( .A(n734), .B(n736), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[9][3] ) );
  INV0 U1167 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[6][5] ), .Q(
        n704) );
  NAND23 U1168 ( .A(n1519), .B(n690), .Q(n1811) );
  XOR30 U1169 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][2] ), .C(n693), .Q(
        n1734) );
  NAND22 U1170 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[4][5] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[5] ), .Q(n1846) );
  XOR22 U1171 ( .A(n1420), .B(n646), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][2] ) );
  INV3 U1172 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[5] ), .Q(n684) );
  XNR31 U1173 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_18_net_[4] ), .B(
        n1518), .C(n707), .Q(n1519) );
  NOR20 U1174 ( .A(n128), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[3] ) );
  INV2 U1175 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[3] ), .Q(n879) );
  INV3 U1176 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[5] ), .Q(
        n1926) );
  NOR20 U1177 ( .A(n128), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[3] ) );
  MAJ32 U1178 ( .A(n1727), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[4] ), .C(n1020), .Q(
        n1520) );
  XOR22 U1179 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[1] ), .Q(n1521) );
  XOR22 U1180 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][1] ), .Q(n1522) );
  NOR21 U1181 ( .A(n145), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[0] ) );
  NOR20 U1182 ( .A(n147), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[4] ) );
  NOR20 U1183 ( .A(n131), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[3] ) );
  INV3 U1184 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[1] ), .Q(n1852) );
  NOR21 U1185 ( .A(n206), .B(n153), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[1] ) );
  INV3 U1186 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[3] ), .Q(n856) );
  INV3 U1187 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_12_net_[3] ), .Q(n477) );
  MAJ31 U1188 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[1][6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[6] ), .C(n589), .Q(n1526) );
  INV3 U1189 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[8][3] ), .Q(
        n547) );
  MAJ31 U1190 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[6] ), .C(n612), .Q(n1527) );
  CLKIN3 U1191 ( .A(n1804), .Q(n1059) );
  XOR21 U1192 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][8] ), .Q(n1528) );
  INV3 U1193 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[1] ), .Q(
        n1929) );
  INV3 U1194 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[1] ), .Q(
        n1732) );
  NOR21 U1195 ( .A(n153), .B(n210), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[1] ) );
  NAND26 U1196 ( .A(n1885), .B(n1884), .Q(n982) );
  NOR21 U1197 ( .A(n131), .B(n203), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[3] ) );
  XNR21 U1198 ( .A(n1594), .B(n410), .Q(n1529) );
  XOR21 U1199 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[3][5] ), .B(
        n638), .Q(n640) );
  IMAJ31 U1200 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[7][4] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[4] ), .C(n1101), .Q(
        n1530) );
  NOR21 U1201 ( .A(n202), .B(n166), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[1] ) );
  NOR23 U1202 ( .A(n148), .B(n193), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[2] ) );
  NAND23 U1203 ( .A(n1849), .B(n1850), .Q(n521) );
  INV3 U1204 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_12_net_[3] ), .Q(n667) );
  INV3 U1205 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[5] ), .Q(
        n1868) );
  XNR21 U1206 ( .A(n1651), .B(n509), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[6][0] ) );
  XNR21 U1207 ( .A(n885), .B(n888), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[6][0] ) );
  INV3 U1208 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[0] ), .Q(
        n1076) );
  INV8 U1209 ( .A(\i_fifo_rx/n154 ), .Q(n302) );
  INV3 U1210 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[2][0] ), .Q(
        n437) );
  INV3 U1211 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[1] ), .Q(n981)
         );
  NAND22 U1212 ( .A(n1915), .B(\i_iq_demod/filtre_Q/out_factor1 [0]), .Q(n1658) );
  NOR21 U1213 ( .A(n200), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[1] ) );
  NOR21 U1214 ( .A(n200), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[1] ) );
  INV3 U1215 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[3] ), .Q(n690) );
  INV8 U1216 ( .A(n1418), .Q(\i_fifo_tx/n6 ) );
  INV8 U1217 ( .A(n1414), .Q(\i_fifo_tx/n7 ) );
  INV8 U1218 ( .A(n1410), .Q(\i_fifo_tx/n8 ) );
  INV8 U1219 ( .A(n1408), .Q(\i_fifo_tx/n9 ) );
  INV8 U1220 ( .A(n1406), .Q(\i_fifo_tx/n73 ) );
  INV8 U1221 ( .A(n124), .Q(\i_fifo_tx/n3 ) );
  INV8 U1222 ( .A(n114), .Q(\i_fifo_tx/n4 ) );
  INV8 U1223 ( .A(n1417), .Q(\i_fifo_rx/n6 ) );
  INV8 U1224 ( .A(n1413), .Q(\i_fifo_rx/n7 ) );
  INV8 U1225 ( .A(n1409), .Q(\i_fifo_rx/n8 ) );
  INV8 U1226 ( .A(n1407), .Q(\i_fifo_rx/n9 ) );
  INV8 U1227 ( .A(n1405), .Q(\i_fifo_rx/n10 ) );
  INV8 U1228 ( .A(n118), .Q(\i_fifo_rx/n4 ) );
  INV8 U1229 ( .A(n112), .Q(\i_fifo_rx/n3 ) );
  INV8 U1230 ( .A(n106), .Q(\i_fifo_rx/n5 ) );
  INV12 U1231 ( .A(n267), .Q(n268) );
  INV12 U1232 ( .A(n265), .Q(n266) );
  BUF12 U1233 ( .A(\i_fifo_rx/N40 ), .Q(n311) );
  INV3 U1234 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[1] ), .Q(
        n1688) );
  NOR21 U1235 ( .A(n153), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[1] ) );
  INV3 U1236 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[3] ), .Q(
        n1866) );
  NOR21 U1237 ( .A(n149), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[1] ) );
  NOR21 U1238 ( .A(n153), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[1] ) );
  INV3 U1239 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_18_net_[1] ), .Q(
        n1613) );
  NOR21 U1240 ( .A(n149), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[1] ) );
  NOR21 U1241 ( .A(n142), .B(n174), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[5] ) );
  NOR21 U1242 ( .A(n156), .B(n166), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[6] ) );
  NOR21 U1243 ( .A(n156), .B(n174), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[6] ) );
  INV3 U1244 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_15_net_[1] ), .Q(
        n1855) );
  NOR21 U1245 ( .A(n202), .B(\i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[1] ) );
  NOR21 U1246 ( .A(n205), .B(n175), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[9] ) );
  NOR21 U1247 ( .A(n166), .B(n212), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[9] ) );
  NOR21 U1248 ( .A(n150), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[4] ) );
  INV3 U1249 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[2] ), .Q(
        n1704) );
  NOR21 U1250 ( .A(n152), .B(n1198), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[2] ) );
  NOR21 U1251 ( .A(n168), .B(n154), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[4] ) );
  INV3 U1252 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_15_net_[3] ), .Q(n500) );
  NOR21 U1253 ( .A(n155), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[6] ) );
  NOR21 U1254 ( .A(n170), .B(n210), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[6] ) );
  NOR21 U1255 ( .A(n199), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[2] ) );
  INV3 U1256 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_15_net_[5] ), .Q(
        n1569) );
  INV3 U1257 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[6] ), .Q(
        n1698) );
  NOR21 U1258 ( .A(n142), .B(\i_iq_demod/filtre_I/mult1_multiplier/n25 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[5] ) );
  NOR21 U1259 ( .A(n199), .B(n1193), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[2] ) );
  NOR31 U1260 ( .A(\i_fifo_rx/n45 ), .B(\i_fifo_rx/n46 ), .C(\i_fifo_rx/n47 ), 
        .Q(\i_fifo_rx/n22 ) );
  NOR31 U1261 ( .A(\i_fifo_tx/n170 ), .B(\i_fifo_tx/n171 ), .C(
        \i_fifo_tx/n172 ), .Q(\i_fifo_tx/n161 ) );
  INV8 U1262 ( .A(n109), .Q(\i_fifo_tx/n5 ) );
  INV3 U1263 ( .A(\i_fifo_rx/n43 ), .Q(\i_fifo_rx/n42 ) );
  INV3 U1264 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[4] ), .Q(
        n1616) );
  INV6 U1265 ( .A(n1568), .Q(n1583) );
  INV3 U1266 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[0] ), .Q(n818)
         );
  NAND22 U1267 ( .A(n1867), .B(n1737), .Q(n1534) );
  CLKIN6 U1268 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][1] ), 
        .Q(n1557) );
  IMAJ30 U1269 ( .A(n1518), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[4] ), .C(n707), .Q(
        n1736) );
  NAND26 U1270 ( .A(n1824), .B(n1825), .Q(n1415) );
  XNR22 U1271 ( .A(n1786), .B(n881), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[6][2] ) );
  XOR31 U1272 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[6][6] ), .C(n890), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[7][5] ) );
  NOR21 U1273 ( .A(n131), .B(n135), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[3] ) );
  XOR21 U1274 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[7] ), .Q(n398) );
  NAND20 U1275 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_9_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][1] ), .Q(n652) );
  NAND26 U1276 ( .A(n1878), .B(n1879), .Q(n1205) );
  XNR22 U1277 ( .A(n1761), .B(n879), .Q(n1668) );
  XOR22 U1278 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[2][7] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[7] ), .Q(n989) );
  AOI221 U1279 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[1][7] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[7] ), .C(n965), .D(
        n966), .Q(n964) );
  NAND23 U1280 ( .A(n1533), .B(n1041), .Q(n1535) );
  NAND22 U1281 ( .A(n1534), .B(n1535), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][4] ) );
  INV3 U1282 ( .A(n1867), .Q(n1533) );
  BUF6 U1283 ( .A(n457), .Q(n1914) );
  MAJ32 U1284 ( .A(n1684), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[4] ), .C(n896), .Q(
        n1536) );
  XNR22 U1285 ( .A(n879), .B(n1761), .Q(n1646) );
  XNR31 U1286 ( .A(n1037), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][6] ), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[6] ), .Q(n1711) );
  NAND22 U1287 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[7][3] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[3] ), .Q(n1789) );
  XNR22 U1288 ( .A(n1705), .B(n1085), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[7][4] ) );
  NAND22 U1289 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[5][5] ), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[5] ), .Q(n1541) );
  NAND26 U1290 ( .A(n1540), .B(n1926), .Q(n1542) );
  NAND28 U1291 ( .A(n1541), .B(n1542), .Q(n875) );
  NAND22 U1292 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][3] ), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[3] ), .Q(n1544) );
  NAND24 U1293 ( .A(n1544), .B(n1545), .Q(n1932) );
  CLKIN3 U1294 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][3] ), 
        .Q(n1543) );
  BUF12 U1295 ( .A(n1932), .Q(n1904) );
  XOR22 U1296 ( .A(n1700), .B(n521), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[7][2] ) );
  XOR21 U1297 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[3][4] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[4] ), .Q(n1546) );
  XOR21 U1298 ( .A(n1720), .B(n1546), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][3] ) );
  XOR22 U1299 ( .A(n1518), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[4] ), .Q(n1547) );
  XOR20 U1300 ( .A(n707), .B(n1547), .Q(n1693) );
  NAND22 U1301 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[4][3] ), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/_12_net_[3] ), .Q(n1875) );
  NOR21 U1302 ( .A(n147), .B(n1187), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[4] ) );
  NAND24 U1303 ( .A(n1615), .B(\i_iq_demod/filtre_Q/out_factor2 [0]), .Q(n1772) );
  IMAJ31 U1304 ( .A(n1684), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[4] ), .C(n896), .Q(
        n1548) );
  NAND22 U1305 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[4][1] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[1] ), .Q(n1550) );
  CLKIN3 U1306 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[4][1] ), 
        .Q(n1549) );
  BUF6 U1307 ( .A(n851), .Q(n1708) );
  XNR22 U1308 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[2] ), .Q(n504) );
  INV2 U1309 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][2] ), .Q(
        net43018) );
  NAND22 U1310 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[6][5] ), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[5] ), .Q(n1859) );
  NAND26 U1311 ( .A(n1564), .B(n879), .Q(n1566) );
  XNR31 U1312 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][8] ), .C(n866), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[6][7] ) );
  INV6 U1313 ( .A(n1679), .Q(n874) );
  NAND21 U1314 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_21_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[7][1] ), .Q(n731) );
  IMAJ31 U1315 ( .A(n727), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[2] ), .C(
        \i_iq_demod/filtre_I/mult2_multiplier/register[7][2] ), .Q(n725) );
  NAND22 U1316 ( .A(n1812), .B(n1553), .Q(n1554) );
  NAND24 U1317 ( .A(n1554), .B(n1555), .Q(n1639) );
  INV2 U1318 ( .A(n1857), .Q(n1553) );
  XOR22 U1319 ( .A(n710), .B(n711), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[7][2] ) );
  INV6 U1320 ( .A(n193), .Q(n1716) );
  INV3 U1321 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[7][3] ), .Q(
        n534) );
  NAND22 U1322 ( .A(n1608), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[4] ), .Q(n1556) );
  AOI220 U1323 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[5][7] ), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[7] ), .C(n1609), .D(
        n868), .Q(n866) );
  XNR20 U1324 ( .A(n553), .B(n555), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[9][0] ) );
  BUF12 U1325 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[6][3] ), .Q(
        n1701) );
  XNR22 U1326 ( .A(n1904), .B(n1667), .Q(n1652) );
  NAND22 U1327 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][1] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[1] ), .Q(n1558) );
  NAND24 U1328 ( .A(n1558), .B(n1559), .Q(n1029) );
  INV3 U1329 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[2] ), .Q(n1560) );
  XOR22 U1330 ( .A(n1934), .B(n1562), .Q(n1933) );
  CLKIN6 U1331 ( .A(n1529), .Q(n1592) );
  XOR31 U1332 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[7][2] ), .C(n1625), .Q(
        n1743) );
  NAND26 U1333 ( .A(n1524), .B(n1877), .Q(n1879) );
  NAND24 U1334 ( .A(n1565), .B(n1566), .Q(n915) );
  XOR31 U1335 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[5][4] ), .B(
        n687), .C(n1616), .Q(n1563) );
  INV6 U1336 ( .A(n1918), .Q(n1002) );
  INV12 U1337 ( .A(n1765), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[1] ) );
  INV6 U1338 ( .A(n1798), .Q(n668) );
  NAND22 U1339 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[7][3] ), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[3] ), .Q(n1565) );
  OAI222 U1340 ( .A(n493), .B(n1569), .C(net41398), .D(n496), .Q(n1568) );
  OAI222 U1341 ( .A(net42042), .B(n1569), .C(net41766), .D(n530), .Q(n528) );
  NAND24 U1342 ( .A(n1571), .B(n1572), .Q(n1570) );
  NAND24 U1343 ( .A(n1575), .B(n1574), .Q(n1573) );
  OAI212 U1344 ( .A(n1583), .B(n1580), .C(n1587), .Q(n1575) );
  CLKIN6 U1345 ( .A(n1573), .Q(n1585) );
  XOR22 U1346 ( .A(n1570), .B(n1586), .Q(n1579) );
  XNR22 U1347 ( .A(n1582), .B(n1583), .Q(n1589) );
  NAND22 U1348 ( .A(n1579), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[5] ), .Q(net41794) );
  BUF2 U1349 ( .A(n433), .Q(net42841) );
  XNR22 U1350 ( .A(n1592), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[2] ), .Q(net43436) );
  IMAJ31 U1351 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_0_net_[3] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[2] ), .C(n411), .Q(n1594) );
  NOR21 U1352 ( .A(n201), .B(n166), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[2] ) );
  OAI312 U1353 ( .A(n1595), .B(n1591), .C(n1590), .D(
        \i_iq_demod/filtre_I/sum1_adder/n14 ), .Q(n1596) );
  OAI311 U1354 ( .A(n1595), .B(n1591), .C(n1590), .D(
        \i_iq_demod/filtre_I/sum1_adder/n14 ), .Q(
        \i_iq_demod/filtre_I/sum1_adder/n8 ) );
  BUF6 U1355 ( .A(net42210), .Q(n1591) );
  XOR21 U1356 ( .A(\i_iq_demod/filtre_I/sum1_adder/n15 ), .B(n1591), .Q(
        net42978) );
  BUF2 U1357 ( .A(n198), .Q(n1595) );
  OAI312 U1358 ( .A(n437), .B(n439), .C(n438), .D(net42565), .Q(n435) );
  BUF4 U1359 ( .A(n435), .Q(net43044) );
  XNR31 U1360 ( .A(n528), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[6] ), .C(
        \i_iq_demod/filtre_I/mult1_multiplier/register[7][6] ), .Q(net41570)
         );
  INV3 U1361 ( .A(net42041), .Q(net42042) );
  INV2 U1362 ( .A(n529), .Q(net42041) );
  NAND24 U1363 ( .A(n529), .B(n1569), .Q(n1597) );
  IMAJ31 U1364 ( .A(n1455), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[4] ), .C(n532), .Q(n530) );
  XOR21 U1365 ( .A(n530), .B(net41766), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[8][4] ) );
  NAND24 U1366 ( .A(net41794), .B(n1597), .Q(net41766) );
  XOR31 U1367 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_12_net_[6] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][6] ), .C(n468), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[5][5] ) );
  INV0 U1368 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][5] ), .Q(
        n493) );
  CLKIN3 U1369 ( .A(net42883), .Q(n1602) );
  OAI222 U1370 ( .A(n470), .B(n471), .C(n472), .D(n473), .Q(n468) );
  XOR22 U1371 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][5] ), .B(
        n471), .Q(n473) );
  CLKIN6 U1372 ( .A(n1598), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][5] ) );
  XNR22 U1373 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_12_net_[5] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][5] ), .Q(n1599) );
  CLKIN1 U1374 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][5] ), 
        .Q(n470) );
  XNR31 U1375 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_9_net_[6] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][6] ), .C(n446), .Q(
        n1598) );
  MAJ32 U1376 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_12_net_[4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][4] ), .C(n474), .Q(
        n1603) );
  OAI222 U1377 ( .A(n1601), .B(n477), .C(n478), .D(net41781), .Q(n474) );
  INV6 U1378 ( .A(n1604), .Q(n478) );
  OAI222 U1379 ( .A(n1601), .B(n477), .C(n478), .D(net41781), .Q(net43064) );
  XOR22 U1380 ( .A(net41781), .B(n478), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[5][2] ) );
  MAJ32 U1381 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[2] ), .C(n480), .Q(
        n1604) );
  NAND23 U1382 ( .A(n1600), .B(n477), .Q(net41833) );
  BUF2 U1383 ( .A(n1600), .Q(n1601) );
  MAJ32 U1384 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[4] ), .C(n497), .Q(
        net42230) );
  IMAJ31 U1385 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[2][4] ), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/_6_net_[4] ), .C(n429), .Q(
        n427) );
  OAI222 U1386 ( .A(net41482), .B(n426), .C(n428), .D(n427), .Q(n423) );
  XOR21 U1387 ( .A(n427), .B(n428), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][4] ) );
  XNR21 U1388 ( .A(n1605), .B(n403), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[2][4] ) );
  INV3 U1389 ( .A(n404), .Q(n1605) );
  NOR20 U1390 ( .A(n154), .B(n166), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[4] ) );
  XOR31 U1391 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_6_net_[4] ), .B(n429), .C(n1606), .Q(net43270) );
  CLKIN3 U1392 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_6_net_[3] ), .Q(
        n432) );
  NAND24 U1393 ( .A(n431), .B(n432), .Q(net41535) );
  OAI222 U1394 ( .A(
        \i_iq_demod/filtre_I/mult1_multiplier/genblk1[0].adder/n10 ), .B(n402), 
        .C(n404), .D(n403), .Q(n400) );
  IMAJ30 U1395 ( .A(\i_iq_demod/filtre_I/data_2_1 [2]), .B(
        \i_iq_demod/filtre_I/data_1_1 [2]), .C(
        \i_iq_demod/filtre_I/sum1_adder/n8 ), .Q(
        \i_iq_demod/filtre_I/sum1_adder/n7 ) );
  XOR21 U1396 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[4] ), .Q(n1788) );
  NAND23 U1397 ( .A(\i_iq_demod/filtre_Q/out_factor2 [3]), .B(n1615), .Q(n1837) );
  INV3 U1398 ( .A(n1710), .Q(n824) );
  NAND23 U1399 ( .A(n1016), .B(n1017), .Q(n1803) );
  NOR21 U1400 ( .A(n461), .B(n459), .Q(n463) );
  NOR21 U1401 ( .A(n154), .B(n138), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[4] ) );
  INV2 U1402 ( .A(n1026), .Q(n1742) );
  CLKIN1 U1403 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[3][3] ), 
        .Q(n643) );
  NAND21 U1404 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][1] ), .Q(n1031) );
  XNR21 U1405 ( .A(n1922), .B(n796), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][0] ) );
  INV6 U1406 ( .A(n1650), .Q(n455) );
  BUF2 U1407 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[5][4] ), .Q(
        n1626) );
  XNR30 U1408 ( .A(n1767), .B(\i_iq_demod/filtre_Q/data_2_2 [2]), .C(
        \i_iq_demod/filtre_Q/data_1_2 [2]), .Q(n204) );
  XOR30 U1409 ( .A(n1614), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[8][2] ), .C(
        \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[2] ), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[9][1] ) );
  BUF2 U1410 ( .A(n1711), .Q(n1813) );
  MAJ32 U1411 ( .A(n1676), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[6] ), .C(net42857), .Q(
        n1748) );
  XOR20 U1412 ( .A(n1867), .B(n1041), .Q(n1610) );
  XOR21 U1413 ( .A(n1522), .B(n842), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][0] ) );
  INV3 U1414 ( .A(n1703), .Q(n1779) );
  XOR22 U1415 ( .A(n1613), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[6][1] ), .Q(n715) );
  BUF2 U1416 ( .A(n740), .Q(n1614) );
  BUF6 U1417 ( .A(n971), .Q(n1686) );
  NAND20 U1418 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[8][1] ), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/_24_net_[1] ), .Q(n744) );
  XOR31 U1419 ( .A(n687), .B(n1685), .C(n1616), .Q(n1712) );
  AOI221 U1420 ( .A(\i_iq_demod/filtre_Q/data_2_2 [3]), .B(
        \i_iq_demod/filtre_Q/data_1_2 [3]), .C(n1218), .D(n1219), .Q(n1217) );
  XOR31 U1421 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[5] ), .B(
        n1617), .C(n1618), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[9][4] ) );
  IMAJ31 U1422 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[8][4] ), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[4] ), .C(n923), .Q(
        n1617) );
  NAND21 U1423 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][1] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[1] ), .Q(n1077) );
  XOR22 U1424 ( .A(n896), .B(n1619), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[7][3] ) );
  BUF2 U1425 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[3][7] ), .Q(
        n1621) );
  XNR22 U1426 ( .A(net42841), .B(net43481), .Q(n1627) );
  AOI221 U1427 ( .A(n1740), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[7] ), .C(n1692), .D(n800), .Q(n798) );
  BUF2 U1428 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[2][6] ), .Q(
        n1622) );
  XNR20 U1429 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[8][3] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[3] ), .Q(n1623) );
  OAI312 U1430 ( .A(n714), .B(n715), .C(n697), .D(n716), .Q(n1624) );
  OAI312 U1431 ( .A(n918), .B(n919), .C(n886), .D(n920), .Q(n1625) );
  OAI311 U1432 ( .A(n919), .B(n918), .C(n886), .D(n920), .Q(n916) );
  XOR22 U1433 ( .A(n1453), .B(n679), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[6][6] ) );
  NAND21 U1434 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][1] ), .Q(n1054) );
  MAJ32 U1435 ( .A(n1648), .B(n1616), .C(n1842), .Q(n720) );
  BUF2 U1436 ( .A(net42078), .Q(net42536) );
  MAJ31 U1437 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[1][7] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[9] ), .C(n396), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[2][8] ) );
  XNR22 U1438 ( .A(net43044), .B(net43436), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][1] ) );
  AOI220 U1439 ( .A(n1696), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[7] ), .C(n1827), .D(n634), .Q(n1628) );
  AOI222 U1440 ( .A(n1740), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[7] ), .C(n1692), .D(n800), .Q(n1629) );
  MAJ32 U1441 ( .A(n1685), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[4] ), .C(n687), .Q(
        n1630) );
  CLKIN3 U1442 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[6][0] ), 
        .Q(n903) );
  XOR22 U1443 ( .A(n852), .B(n1708), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][4] ) );
  IMAJ30 U1444 ( .A(n1614), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[2] ), .C(
        \i_iq_demod/filtre_I/mult2_multiplier/register[8][2] ), .Q(n1631) );
  NOR22 U1445 ( .A(n127), .B(n1892), .Q(n1632) );
  NOR20 U1446 ( .A(n127), .B(n1892), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[3] ) );
  NAND26 U1447 ( .A(n795), .B(n1777), .Q(n1937) );
  XNR21 U1448 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_0_net_[6] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[5] ), .Q(n404) );
  NAND21 U1449 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_12_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][1] ), .Q(n485) );
  XNR22 U1450 ( .A(n1633), .B(n502), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[6][2] ) );
  MAJ31 U1451 ( .A(net43019), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[2] ), .C(n503), .Q(
        n1633) );
  XOR21 U1452 ( .A(n874), .B(n1928), .Q(n1684) );
  BUF2 U1453 ( .A(n167), .Q(n1635) );
  XOR21 U1454 ( .A(n1214), .B(n1216), .Q(n1636) );
  NAND28 U1455 ( .A(n1833), .B(n1834), .Q(net42210) );
  OAI311 U1456 ( .A(n792), .B(n1658), .C(n1937), .D(n795), .Q(n1674) );
  NAND21 U1457 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[7][5] ), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[5] ), .Q(n1840) );
  OAI220 U1458 ( .A(n1620), .B(n1637), .C(n1830), .D(n995), .Q(n991) );
  MAJ31 U1459 ( .A(n1622), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[6] ), .C(n991), .Q(n1647) );
  MAJ32 U1460 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[4][4] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[4] ), .C(n664), .Q(
        n1863) );
  INV3 U1461 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[3] ), .Q(
        n1865) );
  NOR21 U1462 ( .A(n151), .B(n1766), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[4] ) );
  XOR21 U1463 ( .A(n1694), .B(n656), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][6] ) );
  XOR20 U1464 ( .A(n664), .B(n665), .Q(n1640) );
  MAJ31 U1465 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][6] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[6] ), .C(n1015), .Q(
        n1699) );
  NAND22 U1466 ( .A(n997), .B(n999), .Q(n1756) );
  OAI312 U1467 ( .A(n981), .B(n1772), .C(n982), .D(n1884), .Q(n1642) );
  INV6 U1468 ( .A(n1851), .Q(n881) );
  MAJ32 U1469 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[4][2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[2] ), .C(n1739), .Q(
        n1644) );
  XNR22 U1470 ( .A(net43117), .B(n466), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[5][6] ) );
  AOI222 U1471 ( .A(n1761), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[3] ), .C(n1721), .D(
        n1646), .Q(n1645) );
  NAND22 U1472 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][5] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[5] ), .Q(n1802) );
  MAJ32 U1473 ( .A(n1627), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[2] ), .C(n457), .Q(n1650) );
  BUF2 U1474 ( .A(n506), .Q(n1651) );
  XOR22 U1475 ( .A(n1741), .B(n599), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][2] ) );
  IMAJ31 U1476 ( .A(n1664), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[2] ), .C(n600), .Q(n1741) );
  BUF2 U1477 ( .A(n1937), .Q(n1922) );
  CLKBU12 U1478 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[3][2] ), 
        .Q(n1726) );
  MAJ32 U1479 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[2] ), .C(n1072), .Q(
        n1654) );
  NAND23 U1480 ( .A(n1925), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[2] ), .Q(n795) );
  CLKIN2 U1481 ( .A(n1898), .Q(n1666) );
  XNR21 U1482 ( .A(n684), .B(n1883), .Q(n1655) );
  XOR31 U1483 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_9_net_[4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][4] ), .C(n451), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][3] ) );
  NAND24 U1484 ( .A(n1689), .B(n1868), .Q(n1847) );
  NAND26 U1485 ( .A(n1846), .B(n1847), .Q(n1867) );
  XOR20 U1486 ( .A(n1548), .B(n1906), .Q(n1656) );
  MAJ32 U1487 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[1][6] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[6] ), .C(n400), .Q(n1657) );
  NOR20 U1488 ( .A(n1892), .B(n211), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[9] ) );
  NOR20 U1489 ( .A(n207), .B(n1892), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[7] ) );
  NOR20 U1490 ( .A(n155), .B(n1892), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[6] ) );
  NOR21 U1491 ( .A(n150), .B(n1892), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[4] ) );
  NAND23 U1492 ( .A(n1735), .B(n1866), .Q(n1790) );
  XOR21 U1493 ( .A(n1701), .B(n1866), .Q(n1670) );
  BUF2 U1494 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[3][2] ), .Q(
        n1691) );
  IMAJ30 U1495 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[7][2] ), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/_21_net_[2] ), .C(n537), .Q(
        n1659) );
  INV3 U1496 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[8][0] ), .Q(
        n1121) );
  NOR20 U1497 ( .A(n206), .B(n152), .Q(n1660) );
  XOR22 U1498 ( .A(n1216), .B(n1214), .Q(n1661) );
  INV3 U1499 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[0] ), .Q(n1030) );
  CLKIN2 U1500 ( .A(net42758), .Q(net43117) );
  XOR22 U1501 ( .A(n811), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][3] ), .Q(n813) );
  NOR21 U1502 ( .A(n127), .B(n1890), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[3] ) );
  CLKIN1 U1503 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[3] ), .Q(
        n811) );
  OAI312 U1504 ( .A(n602), .B(n1669), .C(n1715), .D(n605), .Q(n1912) );
  OAI312 U1505 ( .A(n524), .B(n525), .C(n507), .D(n526), .Q(n522) );
  NAND21 U1506 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][1] ), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/_15_net_[1] ), .Q(n508) );
  OAI310 U1507 ( .A(n931), .B(n932), .C(n886), .D(n933), .Q(n1665) );
  XNR22 U1508 ( .A(n455), .B(n1666), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][2] ) );
  XNR22 U1509 ( .A(n1904), .B(n1667), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][2] ) );
  XOR22 U1510 ( .A(n1742), .B(n1027), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][1] ) );
  XNR22 U1511 ( .A(n899), .B(n1668), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[7][2] ) );
  NOR21 U1512 ( .A(n144), .B(n1890), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[0] ) );
  XNR22 U1513 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_0_net_[2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[1] ), .Q(n1669) );
  NAND23 U1514 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][1] ), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[1] ), .Q(n819) );
  NAND33 U1515 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[7][0] ), 
        .B(n1714), .C(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[0] ), .Q(
        n1787) );
  BUF2 U1516 ( .A(n1689), .Q(n1672) );
  OAI312 U1517 ( .A(n792), .B(n1658), .C(n1937), .D(n795), .Q(n790) );
  XNR22 U1518 ( .A(n1819), .B(n1673), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][1] ) );
  XNR22 U1519 ( .A(n1759), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[2] ), .Q(n1673) );
  XOR22 U1520 ( .A(n1733), .B(n1035), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][6] ) );
  MAJ31 U1521 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[4][6] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[6] ), .C(n1037), .Q(
        n1733) );
  CLKIN1 U1522 ( .A(n1701), .Q(n1088) );
  XOR21 U1523 ( .A(n1527), .B(n610), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][6] ) );
  XNR31 U1524 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][6] ), .C(n870), .Q(
        n1678) );
  XNR22 U1525 ( .A(n846), .B(n845), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][6] ) );
  MAJ32 U1526 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[4] ), .B(
        n1626), .C(n876), .Q(n1679) );
  CLKIN6 U1527 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[6][3] ), 
        .Q(n1760) );
  MAJ32 U1528 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[3][6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[6] ), .C(n636), .Q(n1827) );
  XOR22 U1529 ( .A(n1680), .B(n1049), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][1] ) );
  XOR22 U1530 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[2] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][2] ), .Q(n1680) );
  CLKIN3 U1531 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[7][0] ), 
        .Q(n1108) );
  NOR20 U1532 ( .A(n1076), .B(n1108), .Q(n1111) );
  INV4 U1533 ( .A(n503), .Q(n1681) );
  CLKIN6 U1534 ( .A(n1681), .Q(n1682) );
  INV3 U1535 ( .A(net43018), .Q(net43019) );
  BUF2 U1536 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][7] ), .Q(
        n1683) );
  MAJ32 U1537 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[6] ), .C(n802), .Q(n1692) );
  OAI312 U1538 ( .A(n525), .B(n524), .C(n507), .D(n526), .Q(n1687) );
  CLKIN3 U1539 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_12_net_[1] ), .Q(
        n1778) );
  NOR21 U1540 ( .A(n202), .B(n174), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[1] ) );
  XOR22 U1541 ( .A(n1779), .B(n1688), .Q(n1094) );
  CLKIN1 U1542 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[3][5] ), 
        .Q(n826) );
  XNR31 U1543 ( .A(n1015), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][6] ), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[6] ), .Q(n1689) );
  XOR31 U1544 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[5][4] ), .B(
        n687), .C(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[4] ), .Q(
        n1690) );
  XNR30 U1545 ( .A(n608), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][8] ), .C(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[9] ), .Q(n1696) );
  XOR21 U1546 ( .A(n1526), .B(n587), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][6] ) );
  NOR22 U1547 ( .A(n146), .B(n1829), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[0] ) );
  NOR21 U1548 ( .A(n142), .B(net42978), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[5] ) );
  CLKIN1 U1549 ( .A(n1905), .Q(n832) );
  XOR22 U1550 ( .A(n1905), .B(n833), .Q(n1697) );
  NAND22 U1551 ( .A(n1711), .B(n1063), .Q(n1887) );
  CLKIN6 U1552 ( .A(n1751), .Q(n834) );
  BUF2 U1553 ( .A(n520), .Q(n1700) );
  XOR31 U1554 ( .A(n1704), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][2] ), .C(n1072), .Q(
        n1703) );
  CLKIN0 U1555 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][5] ), 
        .Q(n849) );
  MAJ32 U1556 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[6][2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[2] ), .C(n712), .Q(
        n1706) );
  CLKIN0 U1557 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[5][3] ), 
        .Q(n878) );
  XOR22 U1558 ( .A(net42210), .B(\i_iq_demod/filtre_I/sum1_adder/n15 ), .Q(
        n1709) );
  MAJ32 U1559 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[3][6] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[6] ), .C(n825), .Q(n1710) );
  CLKIN3 U1560 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_9_net_[0] ), .Q(
        n651) );
  XOR21 U1561 ( .A(n1105), .B(n1104), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[8][2] ) );
  IMAJ31 U1562 ( .A(n1106), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[2] ), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[7][2] ), .Q(n1104) );
  MAJ32 U1563 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][4] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[4] ), .C(n618), .Q(n1713) );
  XOR22 U1564 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[7][1] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[1] ), .Q(n1714) );
  XNR21 U1565 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_0_net_[6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[5] ), .Q(n593) );
  XNR22 U1566 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_0_net_[2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[1] ), .Q(n603) );
  BUF6 U1567 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[8][1] ), .Q(
        n1717) );
  NAND22 U1568 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[8][1] ), .Q(n933) );
  BUF15 U1569 ( .A(n423), .Q(net42857) );
  NOR21 U1570 ( .A(n1008), .B(n1006), .Q(n1010) );
  NAND22 U1571 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_18_net_[1] ), .B(
        n1734), .Q(n716) );
  MAJ32 U1572 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[7][2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[2] ), .C(n916), .Q(
        n1719) );
  XOR22 U1573 ( .A(n691), .B(n692), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[6][2] ) );
  INV6 U1574 ( .A(n1768), .Q(n691) );
  XOR22 U1575 ( .A(n616), .B(n617), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][4] ) );
  NAND21 U1576 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_3_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[2] ), .Q(n605) );
  AOI222 U1577 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][7] ), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/_12_net_[7] ), .C(net42758), 
        .D(n466), .Q(n464) );
  XOR21 U1578 ( .A(n623), .B(n624), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][2] ) );
  MAJ32 U1579 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[6][2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_18_net_[2] ), .C(n901), .Q(
        n1721) );
  XNR30 U1580 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[9] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][8] ), .C(n798), .Q(
        n1722) );
  BUF2 U1581 ( .A(n548), .Q(n1723) );
  XOR22 U1582 ( .A(n450), .B(n449), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][4] ) );
  CLKIN6 U1583 ( .A(n1750), .Q(n449) );
  NAND23 U1584 ( .A(n547), .B(n1930), .Q(n1809) );
  XOR22 U1585 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[8][1] ), .B(
        n1613), .Q(n743) );
  OAI222 U1586 ( .A(n962), .B(n970), .C(n972), .D(n971), .Q(n968) );
  XNR21 U1587 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[6] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[5] ), .Q(n972) );
  XOR21 U1588 ( .A(n1659), .B(n536), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[8][2] ) );
  XNR20 U1589 ( .A(n1059), .B(n1058), .Q(n1730) );
  XNR22 U1590 ( .A(n1731), .B(n1025), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][2] ) );
  INV2 U1591 ( .A(n967), .Q(n965) );
  IMAJ31 U1592 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[1][6] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[6] ), .C(n968), .Q(
        n967) );
  XNR31 U1593 ( .A(n1086), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[6][4] ), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[4] ), .Q(n1735) );
  CLKIN1 U1594 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[8][3] ), 
        .Q(n926) );
  IMAJ31 U1595 ( .A(n1622), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[6] ), .C(n991), .Q(n990)
         );
  XNR21 U1596 ( .A(n967), .B(n966), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][6] ) );
  MAJ32 U1597 ( .A(n1531), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[4] ), .C(n1043), .Q(
        n1737) );
  BUF2 U1598 ( .A(n1119), .Q(n1738) );
  CLKIN3 U1599 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[0] ), .Q(
        n1053) );
  IMAJ31 U1600 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[4] ), .B(
        n1610), .C(n1066), .Q(n1064) );
  BUF2 U1601 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][7] ), .Q(
        n1740) );
  XOR21 U1602 ( .A(n806), .B(n807), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][4] ) );
  IMAJ30 U1603 ( .A(n1663), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[2] ), .C(n1738), .Q(
        n1746) );
  CLKIN1 U1604 ( .A(n1854), .Q(n499) );
  BUF2 U1605 ( .A(n923), .Q(n1747) );
  OAI221 U1606 ( .A(n719), .B(n684), .C(n720), .D(n721), .Q(n718) );
  NOR21 U1607 ( .A(n200), .B(n173), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[1] ) );
  MAJ32 U1608 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[3][4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[4] ), .C(n451), .Q(n1750) );
  MAJ32 U1609 ( .A(n1691), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[2] ), .C(n836), .Q(n1751) );
  NAND22 U1610 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[2][3] ), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/_6_net_[3] ), .Q(n1908) );
  XOR31 U1611 ( .A(n684), .B(n1752), .C(
        \i_iq_demod/filtre_I/mult2_multiplier/register[8][5] ), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[9][4] ) );
  IMAJ31 U1612 ( .A(n734), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[4] ), .C(
        \i_iq_demod/filtre_I/mult2_multiplier/register[8][4] ), .Q(n1752) );
  XOR31 U1613 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[4] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][4] ), .C(n808), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][3] ) );
  CLKIN2 U1614 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_6_net_[3] ), .Q(
        n622) );
  XNR20 U1615 ( .A(n438), .B(n441), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][0] ) );
  CLKIN6 U1616 ( .A(n999), .Q(n1755) );
  NAND22 U1617 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][3] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[3] ), .Q(n1796) );
  INV3 U1618 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][2] ), .Q(
        n1758) );
  INV6 U1619 ( .A(n1758), .Q(n1759) );
  NOR22 U1620 ( .A(n1715), .B(n602), .Q(n606) );
  XOR22 U1621 ( .A(n1745), .B(n1763), .Q(n1762) );
  NAND28 U1622 ( .A(n1415), .B(\i_iq_demod/filtre_I/out_factor2 [1]), .Q(n1765) );
  INV0 U1623 ( .A(n1202), .Q(n1200) );
  NAND22 U1624 ( .A(\i_iq_demod/filtre_I/data_1_2 [1]), .B(n1874), .Q(n1206)
         );
  AOI222 U1625 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[1][7] ), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/_3_net_[7] ), .C(n1657), .D(
        n398), .Q(n396) );
  AOI222 U1626 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[2][7] ), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/_6_net_[7] ), .C(n1748), .D(
        n421), .Q(n419) );
  XOR22 U1627 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[2][7] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[7] ), .Q(n421) );
  XNR21 U1628 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[6][2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[2] ), .Q(n523) );
  BUF6 U1629 ( .A(n1221), .Q(n1767) );
  XNR22 U1630 ( .A(n1726), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[2] ), .Q(n648) );
  NOR21 U1631 ( .A(n140), .B(n1892), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[5] ) );
  NAND26 U1632 ( .A(n1791), .B(n1792), .Q(n1794) );
  CLKIN6 U1633 ( .A(\i_iq_demod/filtre_Q/data_2_2 [1]), .Q(n1791) );
  XOR22 U1634 ( .A(n1862), .B(\i_iq_demod/filtre_Q/data_2_2 [0]), .Q(n1771) );
  XOR22 U1635 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[4][6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[6] ), .Q(n1773) );
  XOR22 U1636 ( .A(n658), .B(n1773), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][5] ) );
  CLKIN6 U1637 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[5][5] ), 
        .Q(n683) );
  NAND22 U1638 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[5][5] ), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[5] ), .Q(n1806) );
  MAJ31 U1639 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][4] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[4] ), .C(n808), .Q(n1889) );
  XNR22 U1640 ( .A(n1419), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[2] ), .Q(n860) );
  XNR22 U1641 ( .A(n1676), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_6_net_[6] ), .Q(n424) );
  INV3 U1642 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[2] ), .Q(n1775) );
  XNR31 U1643 ( .A(n1767), .B(\i_iq_demod/filtre_Q/data_2_2 [2]), .C(
        \i_iq_demod/filtre_Q/data_1_2 [2]), .Q(n1774) );
  OAI310 U1644 ( .A(n197), .B(n163), .C(n1223), .D(n1224), .Q(n1221) );
  INV6 U1645 ( .A(n1925), .Q(n1776) );
  XNR22 U1646 ( .A(net42857), .B(n424), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][5] ) );
  XNR21 U1647 ( .A(n904), .B(n906), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[7][0] ) );
  NOR21 U1648 ( .A(n144), .B(n173), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[0] ) );
  XOR22 U1649 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[5][3] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[3] ), .Q(n1851) );
  XOR22 U1650 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][1] ), .B(
        n1778), .Q(n483) );
  XNR21 U1651 ( .A(n1747), .B(n925), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[9][3] ) );
  XNR21 U1652 ( .A(n1607), .B(n1032), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[4][0] ) );
  IMAJ31 U1653 ( .A(n1707), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[4] ), .C(n853), .Q(n851) );
  NAND22 U1654 ( .A(\i_iq_demod/filtre_Q/data_1_1 [1]), .B(
        \i_iq_demod/filtre_Q/data_2_1 [1]), .Q(n1782) );
  NAND26 U1655 ( .A(n1780), .B(n1781), .Q(n1783) );
  NAND28 U1656 ( .A(n1782), .B(n1783), .Q(n1214) );
  CLKIN6 U1657 ( .A(\i_iq_demod/filtre_Q/data_2_1 [1]), .Q(n1780) );
  CLKIN6 U1658 ( .A(\i_iq_demod/filtre_Q/data_1_1 [1]), .Q(n1781) );
  CLKIN0 U1659 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][5] ), 
        .Q(n804) );
  IMAJ31 U1660 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][6] ), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[6] ), .C(n847), .Q(
        n846) );
  XOR22 U1661 ( .A(n1882), .B(\i_iq_demod/filtre_I/data_2_2 [0]), .Q(n1784) );
  NAND22 U1662 ( .A(\i_iq_demod/filtre_Q/data_1_2 [1]), .B(
        \i_iq_demod/filtre_Q/data_2_2 [1]), .Q(n1793) );
  XOR22 U1663 ( .A(n1785), .B(n1624), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[7][1] ) );
  XOR22 U1664 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_18_net_[2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[6][2] ), .Q(n1785) );
  CLKIN2 U1665 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[3] ), .Q(
        n1001) );
  MAJ32 U1666 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[2] ), .B(
        n1652), .C(n882), .Q(n1786) );
  XOR22 U1667 ( .A(n720), .B(n721), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[8][4] ) );
  XNR22 U1668 ( .A(n1627), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[2] ), .Q(n458) );
  NOR21 U1669 ( .A(n415), .B(n413), .Q(n417) );
  XOR22 U1670 ( .A(n1788), .B(net43064), .Q(n1854) );
  NAND24 U1671 ( .A(n1789), .B(n1790), .Q(n1105) );
  NAND28 U1672 ( .A(n1793), .B(n1794), .Q(n1223) );
  CLKIN6 U1673 ( .A(\i_iq_demod/filtre_Q/data_1_2 [1]), .Q(n1792) );
  INV2 U1674 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[3] ), .Q(n1799) );
  XOR22 U1675 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[8][1] ), .B(
        n1688), .Q(n1122) );
  MAJ32 U1676 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[4][2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[2] ), .C(n670), .Q(
        n1798) );
  INV2 U1677 ( .A(n846), .Q(n844) );
  MAJ31 U1678 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[3][4] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[4] ), .C(n641), .Q(n1800) );
  XOR22 U1679 ( .A(n670), .B(n1801), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][1] ) );
  XOR22 U1680 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[4][2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[2] ), .Q(n1801) );
  OAI312 U1681 ( .A(n884), .B(n885), .C(n886), .D(n887), .Q(n882) );
  XNR30 U1682 ( .A(n1020), .B(n1727), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[4] ), .Q(n1805) );
  AOI221 U1683 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][7] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[7] ), .C(n1804), .D(
        n1058), .Q(n1056) );
  INV3 U1684 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[7][0] ), .Q(
        n729) );
  NAND24 U1685 ( .A(n683), .B(n684), .Q(n1807) );
  XOR22 U1686 ( .A(n668), .B(n1911), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][2] ) );
  NOR22 U1687 ( .A(n484), .B(n482), .Q(n486) );
  NAND22 U1688 ( .A(n1693), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_21_net_[3] ), .Q(n1810) );
  NAND24 U1689 ( .A(n1810), .B(n1811), .Q(n726) );
  XNR22 U1690 ( .A(n635), .B(n634), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][6] ) );
  AOI221 U1691 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[1][7] ), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/_3_net_[7] ), .C(n1526), .D(
        n587), .Q(n585) );
  XNR22 U1692 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_9_net_[5] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][5] ), .Q(n450) );
  OAI312 U1693 ( .A(n195), .B(n161), .C(n1205), .D(n1206), .Q(n1203) );
  AOI221 U1694 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][7] ), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[7] ), .C(n844), .D(
        n845), .Q(n843) );
  XNR31 U1695 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_3_net_[4] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_0_net_[5] ), .C(n594), .Q(n1888) );
  NAND22 U1696 ( .A(\i_iq_demod/filtre_I/data_1_1 [1]), .B(
        \i_iq_demod/filtre_I/data_2_1 [1]), .Q(n1833) );
  AOI221 U1697 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[5][7] ), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[7] ), .C(n1453), .D(
        n679), .Q(n677) );
  XOR31 U1698 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_21_net_[6] ), .B(
        n1815), .C(n718), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[8][5] ) );
  XOR31 U1699 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_18_net_[7] ), .B(
        n1897), .C(n700), .Q(n1815) );
  NAND22 U1700 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][1] ), 
        .B(\i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[1] ), .Q(n1817) );
  CLKIN3 U1701 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][1] ), 
        .Q(n1816) );
  OAI312 U1702 ( .A(n816), .B(n818), .C(n1894), .D(n819), .Q(n1819) );
  XNR21 U1703 ( .A(n862), .B(n865), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][0] ) );
  NAND26 U1704 ( .A(n819), .B(n1839), .Q(n1894) );
  INV0 U1705 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_3_net_[3] ), .Q(n408)
         );
  XOR31 U1706 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[5] ), .B(
        n1820), .C(n1821), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[9][4] ) );
  IMAJ31 U1707 ( .A(n1113), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_24_net_[4] ), .C(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[8][4] ), .Q(n1820) );
  XOR22 U1708 ( .A(net41341), .B(\i_iq_demod/filtre_I/data_2_1 [0]), .Q(n1826)
         );
  XOR22 U1709 ( .A(n1063), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[6][5] ), .Q(n1085) );
  XOR22 U1710 ( .A(net42210), .B(\i_iq_demod/filtre_I/sum1_adder/n15 ), .Q(
        n1828) );
  XOR22 U1711 ( .A(net42210), .B(\i_iq_demod/filtre_I/sum1_adder/n15 ), .Q(
        n1829) );
  XOR22 U1712 ( .A(n1637), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][5] ), .Q(n1830) );
  OAI222 U1713 ( .A(n1678), .B(n873), .C(n1906), .D(n1548), .Q(n890) );
  NAND21 U1714 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][1] ), .Q(n841) );
  NAND26 U1715 ( .A(n1831), .B(n1832), .Q(n1834) );
  CLKIN6 U1716 ( .A(\i_iq_demod/filtre_I/data_2_1 [1]), .Q(n1831) );
  CLKIN6 U1717 ( .A(\i_iq_demod/filtre_I/data_1_1 [1]), .Q(n1832) );
  INV0 U1718 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_9_net_[3] ), .Q(n1899) );
  XOR22 U1719 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][7] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[7] ), .Q(n800) );
  XOR22 U1720 ( .A(n480), .B(n1835), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[5][1] ) );
  XOR22 U1721 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][2] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[2] ), .Q(n1835) );
  XNR31 U1722 ( .A(n677), .B(n1836), .C(
        \i_iq_demod/filtre_I/mult2_multiplier/_15_net_[9] ), .Q(n1897) );
  IMAJ30 U1723 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_12_net_[9] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][8] ), .C(n654), .Q(
        n1836) );
  NOR21 U1724 ( .A(n170), .B(n1766), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[6] ) );
  CLKIN3 U1725 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[6][0] ), 
        .Q(n524) );
  BUF2 U1726 ( .A(n1894), .Q(n1893) );
  INV6 U1727 ( .A(n1856), .Q(n995) );
  NOR21 U1728 ( .A(n143), .B(n203), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[0] ) );
  NAND22 U1729 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[6][3] ), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/_24_net_[3] ), .Q(n1849) );
  NAND24 U1730 ( .A(n1848), .B(n1930), .Q(n1850) );
  INV3 U1731 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_18_net_[3] ), .Q(
        n1930) );
  XNR31 U1732 ( .A(n487), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[5][8] ), .C(
        \i_iq_demod/filtre_I/mult1_multiplier/_15_net_[9] ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[6][7] ) );
  NAND21 U1733 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[7][3] ), 
        .B(\i_iq_demod/filtre_I/mult1_multiplier/_24_net_[3] ), .Q(n1870) );
  OAI312 U1734 ( .A(n539), .B(n540), .C(n507), .D(n541), .Q(n537) );
  XNR22 U1735 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[7][1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_21_net_[1] ), .Q(n540) );
  CLKIN3 U1736 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[7][0] ), 
        .Q(n539) );
  XOR22 U1737 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][1] ), .B(
        n1855), .Q(n506) );
  CLKIN3 U1738 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[5][0] ), 
        .Q(n505) );
  MAJ32 U1739 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[2][4] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[4] ), .C(n997), .Q(n1856) );
  XNR22 U1740 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[1] ), .B(
        n1743), .Q(n932) );
  CLKIN2 U1741 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[8][0] ), 
        .Q(n931) );
  MAJ32 U1742 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[8][2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[2] ), .C(n929), .Q(
        n1858) );
  XNR21 U1743 ( .A(n982), .B(n985), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[2][0] ) );
  XNR22 U1744 ( .A(n1717), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[1] ), .Q(n553) );
  CLKIN2 U1745 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[8][0] ), 
        .Q(n552) );
  OAI312 U1746 ( .A(n602), .B(n603), .C(n1715), .D(n605), .Q(n600) );
  OAI312 U1747 ( .A(n1051), .B(n1053), .C(n1052), .D(n1054), .Q(n1049) );
  OAI312 U1748 ( .A(n552), .B(n553), .C(n507), .D(n554), .Q(n550) );
  XOR22 U1749 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[4][3] ), .B(
        n1865), .Q(n1864) );
  NOR21 U1750 ( .A(n629), .B(n627), .Q(n631) );
  XNR21 U1751 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][2] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[2] ), .Q(n626) );
  AOI222 U1752 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[2][7] ), 
        .B(\i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[7] ), .C(n1647), .D(
        n989), .Q(n987) );
  IMAJ31 U1753 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[6][6] ), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/_18_net_[6] ), .C(n701), .Q(
        n700) );
  NAND21 U1754 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][1] ), .Q(n887) );
  XOR22 U1755 ( .A(n1697), .B(n834), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][2] ) );
  INV3 U1756 ( .A(n1873), .Q(n1874) );
  CLKIN6 U1757 ( .A(\i_iq_demod/filtre_I/data_2_2 [1]), .Q(n1877) );
  BUF2 U1758 ( .A(n414), .Q(net41786) );
  XNR21 U1759 ( .A(n1052), .B(n1055), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[5][0] ) );
  NOR21 U1760 ( .A(n1053), .B(n1051), .Q(n1055) );
  IMAJ30 U1761 ( .A(\i_iq_demod/filtre_I/data_2_2 [2]), .B(
        \i_iq_demod/filtre_I/data_1_2 [2]), .C(n1203), .Q(n1202) );
  IMAJ31 U1762 ( .A(n830), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[4] ), .C(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][4] ), .Q(n828) );
  XNR21 U1763 ( .A(n421), .B(n422), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[3][6] ) );
  OAI312 U1764 ( .A(n1121), .B(n1076), .C(n1122), .D(n1123), .Q(n1119) );
  XNR22 U1765 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[6][1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_18_net_[1] ), .Q(n525) );
  XNR22 U1766 ( .A(n1682), .B(n504), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[6][1] ) );
  INV3 U1767 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[5] ), .Q(
        n1063) );
  NOR21 U1768 ( .A(n148), .B(n203), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[2] ) );
  NOR21 U1769 ( .A(n674), .B(n672), .Q(n676) );
  XOR22 U1770 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[4][5] ), .B(
        n661), .Q(n663) );
  CLKIN1 U1771 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_12_net_[5] ), .Q(
        n661) );
  XNR22 U1772 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_12_net_[4] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][4] ), .Q(n665) );
  CLKIN1 U1773 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_9_net_[3] ), .Q(
        n644) );
  XOR22 U1774 ( .A(n701), .B(n1891), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[7][5] ) );
  XOR22 U1775 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[6][6] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_18_net_[6] ), .Q(n1891) );
  NOR24 U1776 ( .A(n201), .B(n138), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[2] ) );
  XOR21 U1777 ( .A(n788), .B(n789), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[2][2] ) );
  NOR24 U1778 ( .A(n202), .B(n1828), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[1] ) );
  OAI312 U1779 ( .A(n505), .B(n507), .C(n506), .D(n508), .Q(n503) );
  XNR22 U1780 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[3] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[8][3] ), .Q(n928) );
  XNR22 U1781 ( .A(n626), .B(n625), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][1] ) );
  XNR22 U1782 ( .A(n647), .B(n648), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][1] ) );
  XNR22 U1783 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_12_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][1] ), .Q(n673) );
  XOR22 U1784 ( .A(n911), .B(n1902), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[8][3] ) );
  OAI312 U1785 ( .A(n742), .B(n743), .C(n697), .D(n744), .Q(n740) );
  CLKIN2 U1786 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[8][0] ), 
        .Q(n742) );
  XNR22 U1787 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[3] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][3] ), .Q(n692) );
  XOR22 U1788 ( .A(n684), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[7][5] ), .Q(n721) );
  XNR31 U1789 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[4] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[5] ), .C(n973), .Q(n1900) );
  XNR22 U1790 ( .A(n901), .B(n902), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[7][1] ) );
  OAI312 U1791 ( .A(n903), .B(n886), .C(n904), .D(n905), .Q(n901) );
  IMAJ31 U1792 ( .A(n1656), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[4] ), .C(n911), .Q(n909) );
  XOR22 U1793 ( .A(n1101), .B(n1901), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[8][3] ) );
  XOR22 U1794 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[7][4] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_21_net_[4] ), .Q(n1901) );
  CLKIN3 U1795 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[0] ), .Q(
        n840) );
  XOR22 U1796 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[3][7] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[7] ), .Q(n444) );
  XOR22 U1797 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][7] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_12_net_[7] ), .Q(n466) );
  NOR21 U1798 ( .A(n205), .B(n149), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[1] ) );
  XOR21 U1799 ( .A(n593), .B(n592), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][4] ) );
  OAI222 U1800 ( .A(n1482), .B(n1866), .C(n1117), .D(n1118), .Q(n1113) );
  XNR22 U1801 ( .A(n836), .B(n837), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][1] ) );
  CLKBU12 U1802 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[3][3] ), 
        .Q(n1905) );
  XNR22 U1803 ( .A(n1914), .B(n458), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[4][1] ) );
  XNR21 U1804 ( .A(n1853), .B(n1010), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][0] ) );
  CLKIN3 U1805 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[5][0] ), 
        .Q(n884) );
  CLKIN6 U1806 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_0_net_[2] ), .Q(
        n1931) );
  CLKIN3 U1807 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_0_net_[4] ), .Q(
        n407) );
  NOR21 U1808 ( .A(n199), .B(n1890), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[2] ) );
  XOR22 U1809 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[3][7] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[7] ), .Q(n823) );
  XOR31 U1810 ( .A(n1569), .B(net41570), .C(n1936), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[9][4] ) );
  CLKIN1 U1811 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_9_net_[5] ), .Q(
        n638) );
  NAND20 U1812 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[4][1] ), .Q(n864) );
  OAI312 U1813 ( .A(n1634), .B(n650), .C(n651), .D(n652), .Q(n647) );
  INV6 U1814 ( .A(n1909), .Q(n852) );
  XOR22 U1815 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][5] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_12_net_[5] ), .Q(n1909) );
  XNR22 U1816 ( .A(n618), .B(n620), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][3] ) );
  XNR21 U1817 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][4] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[4] ), .Q(n620) );
  XOR22 U1818 ( .A(n639), .B(n640), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[4][4] ) );
  XNR21 U1819 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_24_net_[4] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[8][4] ), .Q(n925) );
  NOR21 U1820 ( .A(n153), .B(n1771), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/_0_net_[1] ) );
  NOR21 U1821 ( .A(n202), .B(n138), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_0_net_[1] ) );
  NOR21 U1822 ( .A(n205), .B(n148), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[2] ) );
  NOR21 U1823 ( .A(n148), .B(n209), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[2] ) );
  XOR21 U1824 ( .A(n812), .B(n813), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][2] ) );
  IMAJ31 U1825 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_0_net_[5] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[4] ), .C(n405), .Q(n403)
         );
  XNR30 U1826 ( .A(n400), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/register[1][6] ), .C(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[6] ), .Q(net41482) );
  XOR22 U1827 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[3][5] ), .B(
        n827), .Q(n1913) );
  CLKIN1 U1828 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[5] ), .Q(
        n827) );
  OAI312 U1829 ( .A(n459), .B(n460), .C(n461), .D(n462), .Q(n457) );
  XNR22 U1830 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[2][5] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_6_net_[5] ), .Q(n807) );
  XNR22 U1831 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_15_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][1] ), .Q(n696) );
  XOR22 U1832 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[2][5] ), .B(
        n426), .Q(n428) );
  CLKIN1 U1833 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_6_net_[5] ), .Q(
        n426) );
  XNR22 U1834 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[3][1] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_9_net_[1] ), .Q(n460) );
  OAI222 U1835 ( .A(n1640), .B(n690), .C(n691), .D(n692), .Q(n687) );
  NOR21 U1836 ( .A(n200), .B(n136), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[1] ) );
  XNR21 U1837 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[2] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[3][2] ), .Q(n837) );
  XNR21 U1838 ( .A(n544), .B(n546), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[9][3] ) );
  XNR22 U1839 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/_15_net_[3] ), .B(
        n1854), .Q(n502) );
  INV0 U1840 ( .A(n1211), .Q(n1209) );
  XNR21 U1841 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[8][4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[4] ), .Q(n546) );
  MAJ32 U1842 ( .A(n1744), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_6_net_[2] ), .C(n1004), .Q(
        n1918) );
  XOR31 U1843 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[7] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[6][7] ), .C(n1079), .Q(
        n1919) );
  NOR24 U1844 ( .A(n162), .B(n196), .Q(n1216) );
  NOR24 U1845 ( .A(n1661), .B(n200), .Q(n1925) );
  XNR22 U1846 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_6_net_[3] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[2][3] ), .Q(n624) );
  XNR22 U1847 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[7][1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_21_net_[1] ), .Q(n919) );
  CLKIN3 U1848 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[7][0] ), 
        .Q(n918) );
  OAI312 U1849 ( .A(n1718), .B(n1030), .C(n1029), .D(n1031), .Q(n1026) );
  XOR22 U1850 ( .A(n1002), .B(n1003), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[3][2] ) );
  IMAJ30 U1851 ( .A(n1730), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_18_net_[6] ), .C(n1080), .Q(
        n1079) );
  XNR22 U1852 ( .A(n1080), .B(n1082), .Q(
        \i_iq_demod/filtre_Q/mult2_multiplier/register[7][5] ) );
  XNR22 U1853 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[5][1] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[1] ), .Q(n885) );
  XNR22 U1854 ( .A(n1931), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_3_net_[1] ), .Q(net41344) );
  CLKIN3 U1855 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[4][0] ), 
        .Q(n672) );
  NOR21 U1856 ( .A(n697), .B(n695), .Q(n699) );
  CLKIN3 U1857 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[6][0] ), 
        .Q(n714) );
  NOR24 U1858 ( .A(n164), .B(n198), .Q(\i_iq_demod/filtre_I/sum1_adder/n15 )
         );
  XOR22 U1859 ( .A(n1905), .B(n833), .Q(n1935) );
  CLKIN1 U1860 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_9_net_[3] ), .Q(
        n833) );
  MAJ32 U1861 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[8][4] ), .B(
        \i_iq_demod/filtre_I/mult1_multiplier/_24_net_[4] ), .C(n544), .Q(
        n1936) );
  XOR22 U1862 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_15_net_[7] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][7] ), .Q(n868) );
  AOI222 U1863 ( .A(n1683), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[7] ), .C(n1699), .D(
        n1013), .Q(n1011) );
  XOR22 U1864 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[3][7] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_9_net_[7] ), .Q(n1013) );
  XOR22 U1865 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[4][7] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_12_net_[7] ), .Q(n1035) );
  OAI312 U1866 ( .A(n1006), .B(n1008), .C(n1762), .D(n1009), .Q(n1004) );
  CLKIN3 U1867 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[4][0] ), 
        .Q(n1051) );
  CLKIN3 U1868 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[2][0] ), 
        .Q(n1006) );
  OAI312 U1869 ( .A(n816), .B(n818), .C(n1894), .D(n819), .Q(n814) );
  OAI312 U1870 ( .A(n861), .B(n863), .C(n862), .D(n864), .Q(n859) );
  OAI222 U1871 ( .A(n704), .B(n684), .C(n1736), .D(n1655), .Q(n701) );
  OAI222 U1872 ( .A(n534), .B(n500), .C(n536), .D(n535), .Q(n532) );
  OAI312 U1873 ( .A(n413), .B(n415), .C(n414), .D(n416), .Q(n411) );
  OAI312 U1874 ( .A(n672), .B(n674), .C(n673), .D(n675), .Q(n670) );
  CLKIN3 U1875 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[4][0] ), 
        .Q(n482) );
  CLKIN3 U1876 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register[3][0] ), 
        .Q(n459) );
  OAI312 U1877 ( .A(n931), .B(n932), .C(n886), .D(n933), .Q(n929) );
  INV3 U1878 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register[4][0] ), .Q(
        n861) );
  XOR22 U1879 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[3][7] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_9_net_[7] ), .Q(n634) );
  AOI222 U1880 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][7] ), 
        .B(\i_iq_demod/filtre_I/mult2_multiplier/_6_net_[7] ), .C(n1527), .D(
        n610), .Q(n608) );
  XOR22 U1881 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][7] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_6_net_[7] ), .Q(n610) );
  XOR22 U1882 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[4][7] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_12_net_[7] ), .Q(n656) );
  XNR22 U1883 ( .A(n882), .B(n883), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[6][1] ) );
  XNR22 U1884 ( .A(n664), .B(n665), .Q(
        \i_iq_demod/filtre_I/mult2_multiplier/register[5][3] ) );
  OAI222 U1885 ( .A(n773), .B(n781), .C(n783), .D(n782), .Q(n779) );
  OAI222 U1886 ( .A(n1540), .B(n873), .C(n874), .D(n875), .Q(n870) );
  OAI312 U1887 ( .A(n1093), .B(n1076), .C(n1094), .D(n1095), .Q(n1091) );
  XNR22 U1888 ( .A(n859), .B(n860), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/register[5][1] ) );
  OAI222 U1889 ( .A(n1088), .B(n1866), .C(n1089), .D(n1090), .Q(n1086) );
  OAI222 U1890 ( .A(n1795), .B(n1799), .C(n1457), .D(n1025), .Q(n1020) );
  OAI222 U1891 ( .A(n1672), .B(n1868), .C(n1041), .D(n1867), .Q(n1037) );
  XOR22 U1892 ( .A(\i_iq_demod/filtre_Q/mult2_multiplier/register[5][7] ), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_15_net_[7] ), .Q(n1058) );
  XNR22 U1893 ( .A(n1687), .B(n523), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/register[7][1] ) );
  OAI222 U1894 ( .A(n878), .B(n879), .C(n880), .D(n881), .Q(n876) );
  OAI222 U1895 ( .A(n926), .B(n879), .C(n927), .D(n928), .Q(n923) );
  OAI222 U1896 ( .A(n810), .B(n811), .C(n812), .D(n813), .Q(n808) );
  OAI222 U1897 ( .A(n1900), .B(n1001), .C(n1002), .D(n1003), .Q(n997) );
  OAI222 U1898 ( .A(n643), .B(n644), .C(n1420), .D(n646), .Q(n641) );
  OAI222 U1899 ( .A(n1848), .B(n500), .C(n521), .D(n520), .Q(n517) );
  OAI222 U1900 ( .A(n447), .B(n448), .C(n449), .D(n450), .Q(n446) );
  OAI222 U1901 ( .A(n583), .B(n591), .C(n593), .D(n592), .Q(n589) );
  OAI222 U1902 ( .A(n849), .B(n850), .C(n852), .D(n851), .Q(n847) );
  OAI222 U1903 ( .A(n1016), .B(n1017), .C(n1869), .D(n1749), .Q(n1015) );
  OAI222 U1904 ( .A(n1813), .B(n1063), .C(n1907), .D(n1064), .Q(n1060) );
  CLKIN3 U1905 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[2][0] ), 
        .Q(n627) );
  OAI222 U1906 ( .A(net42536), .B(n1899), .C(n1898), .D(n455), .Q(n451) );
  OAI222 U1907 ( .A(n407), .B(n408), .C(n410), .D(n409), .Q(n405) );
  IMAJ31 U1908 ( .A(n1638), .B(
        \i_iq_demod/filtre_Q/mult2_multiplier/_3_net_[2] ), .C(n1642), .Q(n977) );
  OAI222 U1909 ( .A(n1724), .B(n667), .C(n668), .D(n1911), .Q(n664) );
  OAI222 U1910 ( .A(n621), .B(n622), .C(n624), .D(n623), .Q(n618) );
  OAI222 U1911 ( .A(n1519), .B(n690), .C(n726), .D(n725), .Q(n722) );
  IMAJ31 U1912 ( .A(n1664), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_3_net_[2] ), .C(n600), .Q(n598)
         );
  OAI222 U1913 ( .A(n826), .B(n827), .C(n1913), .D(n828), .Q(n825) );
  IMAJ31 U1914 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/_0_net_[3] ), .B(
        \i_iq_demod/filtre_Q/mult1_multiplier/_3_net_[2] ), .C(n790), .Q(n788)
         );
  OAI222 U1915 ( .A(n737), .B(n690), .C(n739), .D(n738), .Q(n734) );
  XNR22 U1916 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/_9_net_[1] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/register[3][1] ), .Q(n650) );
  XNR22 U1917 ( .A(\i_iq_demod/filtre_I/mult2_multiplier/register[8][3] ), .B(
        \i_iq_demod/filtre_I/mult2_multiplier/_24_net_[3] ), .Q(n739) );
  NOR31 U1918 ( .A(\i_fifo_tx/n180 ), .B(\i_fifo_tx/n181 ), .C(
        \i_fifo_tx/n182 ), .Q(\i_fifo_tx/n162 ) );
  NOR31 U1919 ( .A(\i_fifo_rx/n153 ), .B(\i_fifo_rx/n154 ), .C(
        \i_fifo_rx/n155 ), .Q(\i_fifo_rx/n23 ) );
  INV3 U1920 ( .A(\i_fifo_rx/n34 ), .Q(\i_fifo_rx/n33 ) );
  INV3 U1921 ( .A(\i_fifo_rx/n169 ), .Q(\i_fifo_rx/n168 ) );
  INV3 U1922 ( .A(\i_fifo_rx/n141 ), .Q(\i_fifo_rx/n140 ) );
  INV3 U1923 ( .A(\i_fifo_rx/n113 ), .Q(\i_fifo_rx/n112 ) );
  INV3 U1924 ( .A(\i_fifo_rx/n88 ), .Q(\i_fifo_rx/n87 ) );
  NOR31 U1925 ( .A(\i_fifo_rx/n154 ), .B(n305), .C(\i_fifo_rx/n155 ), .Q(
        \i_fifo_rx/n29 ) );
  NOR31 U1926 ( .A(n318), .B(\i_fifo_tx/N26 ), .C(\i_fifo_tx/n181 ), .Q(
        \i_fifo_tx/n168 ) );
  INV3 U1927 ( .A(\i_fifo_rx/n83 ), .Q(\i_fifo_rx/n82 ) );
  INV3 U1928 ( .A(\i_fifo_rx/n157 ), .Q(\i_fifo_rx/n156 ) );
  INV3 U1929 ( .A(\i_fifo_rx/n147 ), .Q(\i_fifo_rx/n146 ) );
  INV3 U1930 ( .A(\i_fifo_rx/n124 ), .Q(\i_fifo_rx/n123 ) );
  INV3 U1931 ( .A(\i_fifo_rx/n109 ), .Q(\i_fifo_rx/n108 ) );
  INV3 U1932 ( .A(\i_fifo_rx/n77 ), .Q(\i_fifo_rx/n76 ) );
  INV3 U1933 ( .A(\i_fifo_rx/n64 ), .Q(\i_fifo_rx/n63 ) );
  NOR31 U1934 ( .A(n317), .B(\i_fifo_tx/N26 ), .C(\i_fifo_tx/n180 ), .Q(
        \i_fifo_tx/n167 ) );
  NOR31 U1935 ( .A(\i_fifo_rx/n154 ), .B(\i_fifo_rx/N35 ), .C(\i_fifo_rx/n153 ), .Q(\i_fifo_rx/n35 ) );
  INV3 U1936 ( .A(\i_fifo_rx/n28 ), .Q(\i_fifo_rx/n27 ) );
  INV3 U1937 ( .A(\i_fifo_rx/n151 ), .Q(\i_fifo_rx/n150 ) );
  INV3 U1938 ( .A(\i_fifo_rx/n130 ), .Q(\i_fifo_rx/n129 ) );
  INV3 U1939 ( .A(\i_fifo_rx/n107 ), .Q(\i_fifo_rx/n106 ) );
  INV3 U1940 ( .A(\i_fifo_rx/n86 ), .Q(\i_fifo_rx/n85 ) );
  INV3 U1941 ( .A(\i_fifo_rx/n81 ), .Q(\i_fifo_rx/n80 ) );
  INV3 U1942 ( .A(\i_fifo_rx/n60 ), .Q(\i_fifo_rx/n59 ) );
  NOR31 U1943 ( .A(\i_fifo_tx/n181 ), .B(\i_fifo_tx/N26 ), .C(\i_fifo_tx/n180 ), .Q(\i_fifo_tx/n166 ) );
  INV3 U1944 ( .A(\i_fifo_rx/n163 ), .Q(\i_fifo_rx/n162 ) );
  INV3 U1945 ( .A(\i_fifo_rx/n105 ), .Q(\i_fifo_rx/n104 ) );
  INV3 U1946 ( .A(\i_fifo_rx/n134 ), .Q(\i_fifo_rx/n133 ) );
  INV3 U1947 ( .A(\i_fifo_rx/n37 ), .Q(\i_fifo_rx/n36 ) );
  INV3 U1948 ( .A(\i_fifo_rx/n132 ), .Q(\i_fifo_rx/n131 ) );
  INV3 U1949 ( .A(\i_fifo_rx/n96 ), .Q(\i_fifo_rx/n95 ) );
  INV3 U1950 ( .A(\i_fifo_rx/n69 ), .Q(\i_fifo_rx/n68 ) );
  INV3 U1951 ( .A(\i_fifo_rx/n56 ), .Q(\i_fifo_rx/n55 ) );
  NOR31 U1952 ( .A(n305), .B(\i_fifo_rx/N35 ), .C(\i_fifo_rx/n154 ), .Q(
        \i_fifo_rx/n41 ) );
  NOR31 U1953 ( .A(\i_fifo_tx/n181 ), .B(n318), .C(\i_fifo_tx/n182 ), .Q(
        \i_fifo_tx/n164 ) );
  INV3 U1954 ( .A(\i_fifo_rx/n143 ), .Q(\i_fifo_rx/n142 ) );
  INV3 U1955 ( .A(\i_fifo_rx/n159 ), .Q(\i_fifo_rx/n158 ) );
  INV3 U1956 ( .A(\i_fifo_rx/n117 ), .Q(\i_fifo_rx/n116 ) );
  INV3 U1957 ( .A(\i_fifo_rx/n111 ), .Q(\i_fifo_rx/n110 ) );
  INV3 U1958 ( .A(\i_fifo_rx/n98 ), .Q(\i_fifo_rx/n97 ) );
  INV3 U1959 ( .A(\i_fifo_rx/n73 ), .Q(\i_fifo_rx/n72 ) );
  INV3 U1960 ( .A(\i_fifo_rx/n52 ), .Q(\i_fifo_rx/n51 ) );
  NOR31 U1961 ( .A(\i_fifo_tx/n189 ), .B(\i_fifo_tx/n190 ), .C(
        \i_fifo_tx/n191 ), .Q(\i_fifo_tx/n187 ) );
  NOR31 U1962 ( .A(\i_fifo_tx/n171 ), .B(\i_fifo_tx/N29 ), .C(\i_fifo_tx/n170 ), .Q(\i_fifo_tx/n176 ) );
  NOR31 U1963 ( .A(\i_fifo_rx/n46 ), .B(\i_fifo_rx/N38 ), .C(\i_fifo_rx/n45 ), 
        .Q(\i_fifo_rx/n101 ) );
  INV3 U1964 ( .A(\i_mod_iq/fsm_mapping/n53 ), .Q(\i_mod_iq/fsm_mapping/n119 )
         );
  NAND21 U1965 ( .A(\i_mod_iq/fsm_mapping/C_STATE [1]), .B(
        \i_mod_iq/fsm_mapping/n164 ), .Q(\i_mod_iq/fsm_mapping/n53 ) );
  OAI2112 U1966 ( .A(\i_fifo_rx/n174 ), .B(\i_fifo_rx/n175 ), .C(
        \i_fifo_rx/n176 ), .D(fifo_rx_valid_i), .Q(\i_fifo_rx/n170 ) );
  NAND42 U1967 ( .A(fifo_tx_pwrite_i), .B(n48), .C(fifo_tx_pen_i), .D(
        \i_fifo_tx/n184 ), .Q(\i_fifo_tx/n153 ) );
  INV3 U1968 ( .A(fifo_tx_pslv_err_o), .Q(\i_fifo_tx/n184 ) );
  INV3 U1969 ( .A(\i_fifo_rx/n25 ), .Q(\i_fifo_rx/n24 ) );
  INV3 U1970 ( .A(\i_fifo_rx/n167 ), .Q(\i_fifo_rx/n166 ) );
  INV3 U1971 ( .A(\i_fifo_rx/n145 ), .Q(\i_fifo_rx/n144 ) );
  INV3 U1972 ( .A(\i_fifo_rx/n126 ), .Q(\i_fifo_rx/n125 ) );
  INV3 U1973 ( .A(\i_fifo_rx/n90 ), .Q(\i_fifo_rx/n89 ) );
  INV3 U1974 ( .A(\i_fifo_rx/n54 ), .Q(\i_fifo_rx/n53 ) );
  INV3 U1975 ( .A(\i_fifo_rx/n66 ), .Q(\i_fifo_rx/n65 ) );
  NOR31 U1976 ( .A(n302), .B(\i_fifo_rx/N35 ), .C(\i_fifo_rx/n153 ), .Q(
        \i_fifo_rx/n38 ) );
  NOR31 U1977 ( .A(n302), .B(n305), .C(\i_fifo_rx/n155 ), .Q(\i_fifo_rx/n32 )
         );
  NOR31 U1978 ( .A(\i_fifo_rx/n153 ), .B(n302), .C(\i_fifo_rx/n155 ), .Q(
        \i_fifo_rx/n26 ) );
  INV6 U1979 ( .A(\i_fifo_tx/n181 ), .Q(n317) );
  BUF6 U1980 ( .A(\i_fifo_tx/N31 ), .Q(n327) );
  NOR21 U1981 ( .A(N13), .B(N11), .Q(n73) );
  AOI222 U1982 ( .A(\i_iq_demod/filtre_I/current_state [2]), .B(
        \i_iq_demod/filtre_I/n1 ), .C(\i_iq_demod/filtre_I/n7 ), .D(
        \i_iq_demod/filtre_I/current_state [0]), .Q(\i_iq_demod/filtre_I/n9 )
         );
  AOI222 U1983 ( .A(\i_iq_demod/filtre_Q/current_state [2]), .B(n1384), .C(
        n1388), .D(\i_iq_demod/filtre_Q/current_state [0]), .Q(n1389) );
  NOR31 U1984 ( .A(n317), .B(n319), .C(\i_fifo_tx/n182 ), .Q(\i_fifo_tx/n165 )
         );
  INV3 U1985 ( .A(\i_fifo_rx/n31 ), .Q(\i_fifo_rx/n30 ) );
  INV3 U1986 ( .A(\i_fifo_rx/n103 ), .Q(\i_fifo_rx/n102 ) );
  CLKIN1 U1987 ( .A(\i_fifo_rx/n170 ), .Q(\i_fifo_rx/n171 ) );
  INV3 U1988 ( .A(\i_fifo_rx/n122 ), .Q(\i_fifo_rx/n121 ) );
  INV3 U1989 ( .A(\i_fifo_rx/n165 ), .Q(\i_fifo_rx/n164 ) );
  INV3 U1990 ( .A(\i_fifo_rx/n92 ), .Q(\i_fifo_rx/n91 ) );
  INV3 U1991 ( .A(\i_fifo_rx/n79 ), .Q(\i_fifo_rx/n78 ) );
  INV3 U1992 ( .A(\i_fifo_rx/n49 ), .Q(\i_fifo_rx/n48 ) );
  OAI311 U1993 ( .A(\i_mod_iq/fsm_mapping/n164 ), .B(
        \i_mod_iq/fsm_mapping/n59 ), .C(n252), .D(\i_mod_iq/fsm_mapping/n165 ), 
        .Q(\i_mod_iq/fsm_mapping/n44 ) );
  INV3 U1994 ( .A(\i_fifo_rx/n149 ), .Q(\i_fifo_rx/n148 ) );
  INV6 U1995 ( .A(\i_fifo_tx/n181 ), .Q(n316) );
  XNR20 U1996 ( .A(\i_cordic/cor_y_s0[1][0] ), .B(n360), .Q(\i_cordic/S1/N15 )
         );
  NOR20 U1997 ( .A(n360), .B(\i_cordic/cor_y_s0[1][0] ), .Q(n330) );
  INV2 U1998 ( .A(\i_cordic/cor_x_s0[1][1] ), .Q(n360) );
  NAND22 U1999 ( .A(\i_mod_iq/fsm_mapping/n195 ), .B(
        \i_mod_iq/fsm_mapping/n163 ), .Q(\i_mod_iq/fsm_mapping/n80 ) );
  MUX21 U2000 ( .A(\i_cordic/S1/N15 ), .B(\i_cordic/S1/N21 ), .S(
        \i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/cor_y_s0[2][0] ) );
  MUX21 U2001 ( .A(\i_cordic/S1/N16 ), .B(\i_cordic/S1/N22 ), .S(
        \i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/cor_y_s0[2][1] ) );
  MUX21 U2002 ( .A(\i_cordic/S1/N17 ), .B(\i_cordic/S1/N23 ), .S(
        \i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/cor_y_s0[2][2] ) );
  MUX21 U2003 ( .A(\i_cordic/S1/N18 ), .B(\i_cordic/S1/N24 ), .S(
        \i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/cor_y_s0[2][3] ) );
  MUX21 U2004 ( .A(\i_cordic/S1/N19 ), .B(\i_cordic/S1/N25 ), .S(
        \i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/cor_y_s0[2][4] ) );
  MUX21 U2005 ( .A(\i_cordic/S1/N5 ), .B(\i_cordic/S1/N11 ), .S(
        \i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/cor_x_s0[2][2] ) );
  MUX21 U2006 ( .A(\i_cordic/S1/N6 ), .B(\i_cordic/S1/N12 ), .S(
        \i_cordic/cor_y_s0[1][5] ), .Q(\i_cordic/cor_x_s0[2][3] ) );
  NOR21 U2007 ( .A(n237), .B(\i_mod_iq/fsm_mapping/en_10MHz_prev ), .Q(
        \i_mod_iq/fsm_mapping/N259 ) );
  NOR31 U2008 ( .A(n305), .B(\i_fifo_rx/N35 ), .C(n302), .Q(\i_fifo_rx/n44 )
         );
  NOR31 U2009 ( .A(\i_fifo_tx/n180 ), .B(n317), .C(\i_fifo_tx/n182 ), .Q(
        \i_fifo_tx/n163 ) );
  INV3 U2010 ( .A(\i_iq_demod/filtre_I/sel [0]), .Q(
        \i_iq_demod/filtre_I/data_reg1/n36 ) );
  NOR31 U2011 ( .A(\i_iq_demod/filtre_I/sel [1]), .B(n1943), .C(
        \i_iq_demod/filtre_I/sel [0]), .Q(\i_iq_demod/filtre_I/factor/n5 ) );
  NOR22 U2012 ( .A(\i_iq_demod/filtre_I/n4 ), .B(
        \i_iq_demod/filtre_I/current_state [0]), .Q(
        \i_iq_demod/filtre_I/sel [0]) );
  INV3 U2013 ( .A(\i_iq_demod/filtre_Q/sel [0]), .Q(n1347) );
  NOR31 U2014 ( .A(\i_iq_demod/filtre_Q/sel [1]), .B(n1944), .C(
        \i_iq_demod/filtre_Q/sel [0]), .Q(n1264) );
  NOR22 U2015 ( .A(n1386), .B(\i_iq_demod/filtre_Q/current_state [0]), .Q(
        \i_iq_demod/filtre_Q/sel [0]) );
  INV3 U2016 ( .A(\i_fifo_rx/n71 ), .Q(\i_fifo_rx/n70 ) );
  INV3 U2017 ( .A(\i_fifo_rx/n40 ), .Q(\i_fifo_rx/n39 ) );
  INV3 U2018 ( .A(\i_fifo_rx/n137 ), .Q(\i_fifo_rx/n136 ) );
  INV3 U2019 ( .A(\i_fifo_rx/n100 ), .Q(\i_fifo_rx/n99 ) );
  INV3 U2020 ( .A(\i_fifo_rx/n128 ), .Q(\i_fifo_rx/n127 ) );
  INV3 U2021 ( .A(\i_fifo_rx/n58 ), .Q(\i_fifo_rx/n57 ) );
  NAND22 U2022 ( .A(\i_mod_iq/fsm_mapping/C_STATE [1]), .B(
        \i_mod_iq/fsm_mapping/C_STATE [0]), .Q(\i_mod_iq/fsm_mapping/n90 ) );
  NAND23 U2023 ( .A(N10), .B(n32), .Q(n12) );
  NAND22 U2024 ( .A(sel_i[0]), .B(n81), .Q(N10) );
  NOR31 U2025 ( .A(\i_fifo_tx/N28 ), .B(\i_fifo_tx/N29 ), .C(\i_fifo_tx/n171 ), 
        .Q(\i_fifo_tx/n178 ) );
  NOR31 U2026 ( .A(\i_fifo_tx/n171 ), .B(\i_fifo_tx/N28 ), .C(\i_fifo_tx/n172 ), .Q(\i_fifo_tx/n174 ) );
  NOR31 U2027 ( .A(\i_fifo_rx/N37 ), .B(\i_fifo_rx/N38 ), .C(\i_fifo_rx/n46 ), 
        .Q(\i_fifo_rx/n135 ) );
  NOR31 U2028 ( .A(\i_fifo_rx/n46 ), .B(\i_fifo_rx/N37 ), .C(\i_fifo_rx/n47 ), 
        .Q(\i_fifo_rx/n67 ) );
  CLKIN6 U2029 ( .A(\i_fifo_rx/n153 ), .Q(n303) );
  BUF6 U2030 ( .A(\i_fifo_tx/N31 ), .Q(n328) );
  INV6 U2031 ( .A(\i_fifo_tx/n181 ), .Q(n314) );
  INV6 U2032 ( .A(\i_fifo_rx/n154 ), .Q(n300) );
  NOR41 U2033 ( .A(n244), .B(n394), .C(n393), .D(n392), .Q(\i_cdr/i_cdr/N145 )
         );
  INV3 U2034 ( .A(\i_iq_demod/filtre_I/factor/n8 ), .Q(
        \i_iq_demod/filtre_I/factor/n24 ) );
  INV3 U2035 ( .A(n1267), .Q(n1269) );
  INV3 U2036 ( .A(\i_cordic/n19 ), .Q(\i_cordic/cor_x_s0[0][3] ) );
  INV3 U2037 ( .A(\i_cordic/n20 ), .Q(\i_cordic/cor_x_s0[0][2] ) );
  INV3 U2038 ( .A(\i_cordic/n21 ), .Q(\i_cordic/cor_x_s0[0][1] ) );
  XNR21 U2039 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register_pipe[11][1] ), .B(\i_iq_demod/filtre_I/mult1_multiplier/_51_net_[1] ), .Q(n577) );
  XNR21 U2040 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/register_pipe[10][1] ), .B(\i_iq_demod/filtre_I/mult1_multiplier/_51_net_[1] ), .Q(n571) );
  INV3 U2041 ( .A(\i_iq_demod/filtre_I/mult1_multiplier/n20 ), .Q(
        \i_iq_demod/filtre_I/mult1_multiplier/_51_net_[1] ) );
  XNR21 U2042 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[11][1] ), .B(\i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[1] ), .Q(n956) );
  XNR21 U2043 ( .A(\i_iq_demod/filtre_Q/mult1_multiplier/register_pipe[10][1] ), .B(\i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[1] ), .Q(n950) );
  INV3 U2044 ( .A(n1191), .Q(
        \i_iq_demod/filtre_Q/mult1_multiplier/_51_net_[1] ) );
  AOI221 U2045 ( .A(\i_cordic/S2/N20 ), .B(n185), .C(\i_cordic/cor_y_s1[2][5] ), .D(\i_cordic/S2/N26 ), .Q(\i_cordic/S2/n21 ) );
  NOR31 U2046 ( .A(n319), .B(\i_fifo_tx/N26 ), .C(n317), .Q(\i_fifo_tx/n169 )
         );
  NAND22 U2047 ( .A(\i_mod_iq/fsm_mapping/n56 ), .B(\i_mod_iq/fsm_mapping/n57 ), .Q(\i_mod_iq/fsm_mapping/n92 ) );
  CLKIN0 U2048 ( .A(n85), .Q(\i_mod_iq/fsm_mapping/n57 ) );
  INV3 U2049 ( .A(n1938), .Q(n1939) );
  INV3 U2050 ( .A(\i_fifo_rx/n172 ), .Q(\i_fifo_rx/n173 ) );
  INV3 U2051 ( .A(n1940), .Q(n1941) );
  OAI312 U2052 ( .A(\i_cordic/n5 ), .B(\i_cordic/qbb_ibuff [4]), .C(
        \i_cordic/n6 ), .D(\i_cordic/n7 ), .Q(n1942) );
  OAI211 U2053 ( .A(n1942), .B(\i_cordic/S0/n22 ), .C(\i_cordic/S0/n33 ), .Q(
        \i_cordic/cor_x_s0[1][4] ) );
  XNR20 U2054 ( .A(n1942), .B(\i_cordic/S0/r64/carry [5]), .Q(n277) );
  OAI221 U2055 ( .A(\i_cordic/S0/n39 ), .B(\i_cordic/S0/n22 ), .C(n1942), .D(
        \i_cordic/S0/n23 ), .Q(\i_cordic/cor_y_s0[1][4] ) );
  OAI221 U2056 ( .A(\i_cordic/S0/n39 ), .B(\i_cordic/S0/n26 ), .C(n1942), .D(
        \i_cordic/S0/n27 ), .Q(\i_cordic/cor_y_s0[1][2] ) );
  OAI211 U2057 ( .A(n1942), .B(\i_cordic/S0/n24 ), .C(\i_cordic/S0/n34 ), .Q(
        \i_cordic/cor_x_s0[1][3] ) );
  OAI221 U2058 ( .A(\i_cordic/S0/n39 ), .B(\i_cordic/S0/n24 ), .C(n1942), .D(
        \i_cordic/S0/n25 ), .Q(\i_cordic/cor_y_s0[1][3] ) );
  OAI211 U2059 ( .A(n1942), .B(\i_cordic/S0/n26 ), .C(\i_cordic/S0/n35 ), .Q(
        \i_cordic/cor_x_s0[1][2] ) );
  OAI221 U2060 ( .A(\i_cordic/S0/n39 ), .B(\i_cordic/S0/n28 ), .C(n1942), .D(
        \i_cordic/S0/n29 ), .Q(\i_cordic/cor_y_s0[1][1] ) );
  INV3 U2061 ( .A(\i_cordic/cor_y_s0[0][5] ), .Q(\i_cordic/S0/n39 ) );
  OAI311 U2062 ( .A(\i_cordic/n5 ), .B(\i_cordic/qbb_ibuff [4]), .C(
        \i_cordic/n6 ), .D(\i_cordic/n7 ), .Q(\i_cordic/cor_y_s0[0][5] ) );
  NOR21 U2063 ( .A(\i_mod_iq/fsm_mapping/n40 ), .B(\i_mod_iq/fsm_mapping/n127 ), .Q(\i_mod_iq/fsm_mapping/n39 ) );
  NOR21 U2064 ( .A(\i_mod_iq/fsm_mapping/N259 ), .B(
        \i_mod_iq/fsm_mapping/n127 ), .Q(\i_mod_iq/fsm_mapping/n40 ) );
  INV3 U2065 ( .A(\i_fifo_rx/n62 ), .Q(\i_fifo_rx/n61 ) );
  INV3 U2066 ( .A(\i_fifo_rx/n94 ), .Q(\i_fifo_rx/n93 ) );
  INV3 U2067 ( .A(\i_fifo_rx/n75 ), .Q(\i_fifo_rx/n74 ) );
  INV3 U2068 ( .A(\i_fifo_rx/n161 ), .Q(\i_fifo_rx/n160 ) );
  INV3 U2069 ( .A(\i_fifo_rx/n139 ), .Q(\i_fifo_rx/n138 ) );
  INV3 U2070 ( .A(\i_fifo_rx/n120 ), .Q(\i_fifo_rx/n119 ) );
  INV3 U2071 ( .A(\i_fifo_rx/n115 ), .Q(\i_fifo_rx/n114 ) );
  INV3 U2072 ( .A(\i_fifo_rx/n14 ), .Q(\i_fifo_rx/n12 ) );
  NOR22 U2073 ( .A(n49), .B(n5), .Q(n51) );
  INV3 U2074 ( .A(n32), .Q(n49) );
  NAND22 U2075 ( .A(N12), .B(n32), .Q(n4) );
  NAND22 U2076 ( .A(sel_i[1]), .B(n80), .Q(N12) );
  NAND22 U2077 ( .A(\i_iq_demod/sine_IN [1]), .B(\i_iq_demod/sine_IN [0]), .Q(
        \i_iq_demod/demod/n20 ) );
  NAND22 U2078 ( .A(\i_iq_demod/cosine_IN [1]), .B(\i_iq_demod/cosine_IN [0]), 
        .Q(\i_iq_demod/demod/n32 ) );
  NAND22 U2079 ( .A(\i_fifo_tx/state_rd ), .B(\i_fifo_tx/n191 ), .Q(
        \i_fifo_tx/n81 ) );
  NAND30 U2080 ( .A(\i_fifo_tx/counter_clock [4]), .B(
        \i_fifo_tx/counter_clock [3]), .C(\i_fifo_tx/n203 ), .Q(
        \i_fifo_tx/n191 ) );
  CLKIN1 U2081 ( .A(n1311), .Q(n1943) );
  AOI210 U2082 ( .A(\i_iq_demod/filtre_I/data_reg1/n36 ), .B(
        \i_iq_demod/filtre_I/n9 ), .C(n1943), .Q(
        \i_iq_demod/filtre_I/out_factor1_req [3]) );
  IMUX20 U2083 ( .A(n1943), .B(\i_iq_demod/filtre_I/sel [0]), .S(
        \i_iq_demod/filtre_I/n9 ), .Q(\i_iq_demod/filtre_I/out_factor2_req [6]) );
  AOI210 U2084 ( .A(\i_iq_demod/filtre_I/sel [0]), .B(\i_iq_demod/filtre_I/n9 ), .C(n1943), .Q(\i_iq_demod/filtre_I/out_factor2_req [4]) );
  NOR30 U2085 ( .A(\i_iq_demod/filtre_I/sel [1]), .B(n1943), .C(
        \i_iq_demod/filtre_I/data_reg1/n36 ), .Q(
        \i_iq_demod/filtre_I/factor/n4 ) );
  NOR30 U2086 ( .A(\i_iq_demod/filtre_I/data_reg1/n36 ), .B(
        \i_iq_demod/filtre_I/sel [2]), .C(\i_iq_demod/filtre_I/n9 ), .Q(
        \i_iq_demod/filtre_I/factor/n8 ) );
  NOR31 U2087 ( .A(\i_iq_demod/filtre_I/data_reg1/n36 ), .B(
        \i_iq_demod/filtre_I/sel [2]), .C(\i_iq_demod/filtre_I/n9 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n8 ) );
  NOR31 U2088 ( .A(\i_iq_demod/filtre_I/data_reg1/n36 ), .B(
        \i_iq_demod/filtre_I/sel [2]), .C(\i_iq_demod/filtre_I/n9 ), .Q(n1283)
         );
  NOR31 U2089 ( .A(\i_iq_demod/filtre_I/sel [0]), .B(
        \i_iq_demod/filtre_I/sel [2]), .C(\i_iq_demod/filtre_I/n9 ), .Q(
        \i_iq_demod/filtre_I/data_reg1/n6 ) );
  NOR31 U2090 ( .A(\i_iq_demod/filtre_I/sel [0]), .B(
        \i_iq_demod/filtre_I/sel [2]), .C(\i_iq_demod/filtre_I/n9 ), .Q(n1281)
         );
  NOR31 U2091 ( .A(\i_iq_demod/filtre_I/sel [1]), .B(
        \i_iq_demod/filtre_I/sel [2]), .C(\i_iq_demod/filtre_I/sel [0]), .Q(
        \i_iq_demod/filtre_I/data_reg1/n5 ) );
  NOR31 U2092 ( .A(\i_iq_demod/filtre_I/sel [1]), .B(
        \i_iq_demod/filtre_I/sel [2]), .C(\i_iq_demod/filtre_I/sel [0]), .Q(
        n1280) );
  CLKIN1 U2093 ( .A(n1348), .Q(n1944) );
  AOI210 U2094 ( .A(n1347), .B(n1389), .C(n1944), .Q(
        \i_iq_demod/filtre_Q/out_factor1_req [3]) );
  IMUX20 U2095 ( .A(n1944), .B(\i_iq_demod/filtre_Q/sel [0]), .S(n1389), .Q(
        \i_iq_demod/filtre_Q/out_factor2_req [6]) );
  AOI210 U2096 ( .A(\i_iq_demod/filtre_Q/sel [0]), .B(n1389), .C(n1944), .Q(
        \i_iq_demod/filtre_Q/out_factor2_req [4]) );
  NOR30 U2097 ( .A(\i_iq_demod/filtre_Q/sel [1]), .B(n1944), .C(n1347), .Q(
        n1263) );
  NOR30 U2098 ( .A(n1347), .B(\i_iq_demod/filtre_Q/sel [2]), .C(n1389), .Q(
        n1267) );
  NOR31 U2099 ( .A(n1347), .B(\i_iq_demod/filtre_Q/sel [2]), .C(n1389), .Q(
        n1356) );
  NOR31 U2100 ( .A(n1347), .B(\i_iq_demod/filtre_Q/sel [2]), .C(n1389), .Q(
        n1319) );
  NOR31 U2101 ( .A(\i_iq_demod/filtre_Q/sel [0]), .B(
        \i_iq_demod/filtre_Q/sel [2]), .C(n1389), .Q(n1354) );
  NOR31 U2102 ( .A(\i_iq_demod/filtre_Q/sel [0]), .B(
        \i_iq_demod/filtre_Q/sel [2]), .C(n1389), .Q(n1317) );
  NOR31 U2103 ( .A(\i_iq_demod/filtre_Q/sel [1]), .B(
        \i_iq_demod/filtre_Q/sel [2]), .C(\i_iq_demod/filtre_Q/sel [0]), .Q(
        n1353) );
  NOR31 U2104 ( .A(\i_iq_demod/filtre_Q/sel [1]), .B(
        \i_iq_demod/filtre_Q/sel [2]), .C(\i_iq_demod/filtre_Q/sel [0]), .Q(
        n1316) );
  INV3 U2105 ( .A(\i_iq_demod/filtre_Q/sel [2]), .Q(n1348) );
  INV2 U2106 ( .A(\i_mod_iq/fsm_mapping/n68 ), .Q(\i_mod_iq/fsm_mapping/n51 )
         );
  NAND22 U2107 ( .A(\i_mod_iq/fsm_mapping/n68 ), .B(
        \i_mod_iq/fsm_mapping/cpt [2]), .Q(\i_mod_iq/fsm_mapping/n76 ) );
  NOR21 U2108 ( .A(\i_mod_iq/fsm_mapping/n47 ), .B(\i_mod_iq/fsm_mapping/n68 ), 
        .Q(\i_mod_iq/fsm_mapping/n193 ) );
  AOI2111 U2109 ( .A(\i_mod_iq/fsm_mapping/n175 ), .B(
        \i_mod_iq/fsm_mapping/n131 ), .C(\i_mod_iq/fsm_mapping/n127 ), .D(
        \i_mod_iq/fsm_mapping/n68 ), .Q(\i_mod_iq/fsm_mapping/n167 ) );
  NOR21 U2110 ( .A(\i_mod_iq/fsm_mapping/n164 ), .B(
        \i_mod_iq/fsm_mapping/C_STATE [1]), .Q(\i_mod_iq/fsm_mapping/n68 ) );
  INV3 U2111 ( .A(\i_fifo_rx/n155 ), .Q(n1945) );
  INV3 U2112 ( .A(\i_fifo_tx/n182 ), .Q(n1946) );
  INV6 U2113 ( .A(n271), .Q(n272) );
  INV6 U2114 ( .A(n269), .Q(n270) );
  NAND33 U2115 ( .A(n104), .B(n105), .C(\i_fifo_rx/n217 ), .Q(\i_fifo_rx/n188 ) );
  NOR31 U2116 ( .A(\i_fifo_rx/i [5]), .B(\i_fifo_rx/i [7]), .C(
        \i_fifo_rx/i [6]), .Q(\i_fifo_rx/n217 ) );
  NOR31 U2117 ( .A(\i_fifo_tx/N28 ), .B(\i_fifo_tx/N29 ), .C(n273), .Q(
        \i_fifo_tx/n179 ) );
  NOR31 U2118 ( .A(n273), .B(\i_fifo_tx/N28 ), .C(\i_fifo_tx/n172 ), .Q(
        \i_fifo_tx/n175 ) );
  NOR31 U2119 ( .A(n273), .B(\i_fifo_tx/N29 ), .C(\i_fifo_tx/n170 ), .Q(
        \i_fifo_tx/n177 ) );
  NOR31 U2120 ( .A(\i_fifo_tx/n170 ), .B(n273), .C(\i_fifo_tx/n172 ), .Q(
        \i_fifo_tx/n173 ) );
  NOR31 U2121 ( .A(\i_fifo_rx/N37 ), .B(\i_fifo_rx/N38 ), .C(n274), .Q(
        \i_fifo_rx/n152 ) );
  NOR31 U2122 ( .A(n274), .B(\i_fifo_rx/N37 ), .C(\i_fifo_rx/n47 ), .Q(
        \i_fifo_rx/n84 ) );
  NOR31 U2123 ( .A(n274), .B(\i_fifo_rx/N38 ), .C(\i_fifo_rx/n45 ), .Q(
        \i_fifo_rx/n118 ) );
  NOR31 U2124 ( .A(\i_fifo_rx/n45 ), .B(n274), .C(\i_fifo_rx/n47 ), .Q(
        \i_fifo_rx/n50 ) );
  CLKIN6 U2125 ( .A(\i_fifo_tx/n181 ), .Q(n315) );
  CLKIN6 U2126 ( .A(\i_fifo_rx/n154 ), .Q(n299) );
  BUF6 U2127 ( .A(\i_fifo_tx/N31 ), .Q(n326) );
  INV6 U2128 ( .A(\i_fifo_rx/n153 ), .Q(n305) );
  CLKIN1 U2129 ( .A(\i_fifo_tx/n153 ), .Q(\i_fifo_tx/n152 ) );
  INV8 U2130 ( .A(\i_fifo_tx/n180 ), .Q(n319) );
  CLKIN8 U2131 ( .A(\i_fifo_tx/n180 ), .Q(n318) );
  INV12 U2132 ( .A(n133), .Q(n306) );
  INV12 U2133 ( .A(n133), .Q(n307) );
  INV12 U2134 ( .A(n126), .Q(n324) );
  INV12 U2135 ( .A(n126), .Q(n321) );
endmodule

